//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   ICLAB 2023 Fall
//   Lab01 Exercise     : Snack Shopping Calculator
//   Author             : Yu-Hsiang Wang
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : V1.0 (Release Date: 2024-09)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

`define CYCLE_TIME 20.0

`ifdef RTL
    `define PATTERN_NUM 40
`endif
`ifdef GATE
    `define PATTERN_NUM 40
`endif

module PATTERN(
  // Output signals
    card_num,
    input_money,
    snack_num,
    price, 
  // Input signals
    out_valid,
    out_change
);

//================================================================
//   INPUT AND OUTPUT DECLARATION                         
//================================================================
output reg [63:0] card_num;
output reg [8:0] input_money;
output reg [31:0] snack_num;
output reg [31:0] price;
input out_valid;
input [8:0] out_change;

//================================================================
// parameters & integer
//================================================================
integer PATNUM = 10000;
integer patcount;
integer input_file, output_file;
integer k,i,j;

//================================================================
// wire & registers 
//================================================================
reg [3:0] golden_card_num [0:15];
reg [8:0] golden_input_money;
reg [3:0] golden_snack_num [0:7];
reg [3:0] golden_price [0:7];
reg golden_valid;
reg [8:0] golden_change;

//================================================================
// clock
//================================================================
reg clk;
real    CYCLE = `CYCLE_TIME;
always  #(CYCLE/2.0) clk = ~clk;
initial clk = 0;

//================================================================
// Hint
//================================================================
// if you want to use c++/python to generate test data, here is 
// a sample format for you. You can change for your convinience.
/* input.txt format
1. [PATTERN_NUM] 

repeat(PATTERN_NUM)
    1. [card_num_0] [card_num_1] ... [card_num_15} 
    2. [input_money]
    3. [snack_num_0] [snack_num_1] ... [snack_num_7]
    4. [price_0] [price_1] ... [price_7]
*/

/* output.txt format
1. [out_valid]
2. [out_change]
*/

//================================================================
// initial
//================================================================
initial begin
    input_file=$fopen("../00_TESTBED/input.txt","r");
    output_file=$fopen("../00_TESTBED/output.txt","r");

    card_num = 'bx;
    input_money = 'bx;
    snack_num = 'bx;
    price = 'bx;
    repeat(5) @(negedge clk);

    k = $fscanf(input_file, "%d", PATNUM);

    for( patcount = 0; patcount < PATNUM; patcount=patcount+1) begin        
        input_task;
        repeat(1) @(negedge clk);
        check_ans;
        repeat($urandom_range(3, 5)) @(negedge clk);
    end
    display_pass;
    repeat(3) @(negedge clk);
    $finish;
end

//================================================================
// task
//================================================================

task input_task; begin
    // k = $fscanf(input_file,"%d",parameter);
    for ( i = 0; i < 16; i=i+1) begin
        k = $fscanf(input_file, "%d", golden_card_num[i]);
    end

    k = $fscanf(input_file, "%d", golden_input_money);

    for ( i = 0; i < 8; i=i+1) begin
        k = $fscanf(input_file, "%d", golden_snack_num[i]);
    end

    for ( i = 0; i < 8; i=i+1) begin
        k = $fscanf(input_file, "%d", golden_price[i]);
    end

    card_num = {golden_card_num[0], golden_card_num[1], golden_card_num[2], golden_card_num[3], 
                golden_card_num[4], golden_card_num[5], golden_card_num[6], golden_card_num[7], 
                golden_card_num[8], golden_card_num[9], golden_card_num[10], golden_card_num[11], 
                golden_card_num[12], golden_card_num[13], golden_card_num[14], golden_card_num[15]};
    input_money = golden_input_money;
    snack_num = {golden_snack_num[0], golden_snack_num[1], golden_snack_num[2], golden_snack_num[3], 
                 golden_snack_num[4], golden_snack_num[5], golden_snack_num[6], golden_snack_num[7]};
    price = {golden_price[0], golden_price[1], golden_price[2], golden_price[3], 
             golden_price[4], golden_price[5], golden_price[6], golden_price[7]};

end endtask

task check_ans; begin
    // k = $fscanf(output_file,"%d",golden_ans);  
    k = $fscanf(output_file,"%d",golden_valid);
    k = $fscanf(output_file,"%d",golden_change);
    if(out_valid !== golden_valid) begin
        display_fail;
        $display ("-------------------------------------------------------------------");
        $display("*                            PATTERN NO.%4d 	                      ", patcount);
        $display ("         card valid should be : %d , your answer is : %d           ", golden_valid, out_valid);
        $display ("-------------------------------------------------------------------");
        #(100);
        $finish ;
    end
    else if (out_change !== golden_change) begin
        display_fail;
        $display ("-------------------------------------------------------------------");
        $display("*                            PATTERN NO.%4d 	                      ", patcount);
        $display ("            change should be : %d , your answer is : %d           ", golden_change, out_change);
        $display ("-------------------------------------------------------------------");
        #(100);
        $finish ;
    end
    else $display ("             \033[0;32mPass Pattern NO. %d\033[m         ", patcount);
end endtask

task display_fail; begin
    $display("\n");
    $display("\n");
    $display("\033[0;37m....................................................................................................\033[0m");
    $display("\033[0;37m.......................................................................,:+++:.......................\033[0m");
    $display("\033[0;37m....................................................,:+*\033[0m\033[0;32m******\033[0m\033[0;37m+;,....:*\033[0m\033[0;30m%%%%?%%S\033[0m\033[0;37m.\033[0m\033[0;30mS\033[0m\033[0;37m*:....................\033[0m");
    $display("\033[0;37m................................................,:*\033[0m\033[0;30m?%%%%%%%%\033[0m\033[0;32m????\033[0m\033[0;30m?%%%%%%%%\033[0m\033[0;32m*\033[0m\033[0;37m:.;.\033[0m\033[0;30m%%\033[0m\033[0;32m?\033[0m\033[0;30m%%SS%%%%SSS%%\033[0m\033[0;37m:..................\033[0m");
    $display("\033[0;37m..............................................:+\033[0m\033[0;30m?%%%%\033[0m\033[0;32m?????\033[0m\033[0;30m%%SSSSSSSSSSS\033[0m\033[0;37m.\033[0m\033[0;30m%%%%SSSSSS%%%%%%S\033[0m\033[0;37m.*,................\033[0m");
    $display("\033[0;37m...........................................:+\033[0m\033[0;30m?%%%%\033[0m\033[0;32m??????\033[0m\033[0;30mSS%%%%%%%%SSSSS#\033[0m\033[0;37m..\033[0m\033[0;30mSSSSS%%\033[0m\033[0;32m???????\033[0m\033[0;30m%%SS\033[0m\033[0;37m;...............\033[0m");
    $display("\033[0;37m........................................:+\033[0m\033[0;30m?%%%%\033[0m\033[0;32m???????\033[0m\033[0;30m%%S%%?%%SS%%%%???%%%%%%\033[0m\033[0;37m..\033[0m\033[0;30mSS%%\033[0m\033[0;32m??\033[0m\033[0;30m%%%%%%%%?\033[0m\033[0;32m*\033[0m\033[0;37m***\033[0m\033[0;30m?S\033[0m\033[0;37m*..............\033[0m");
    $display("\033[0;37m....................................,:+\033[0m\033[0;30m?%%%%\033[0m\033[0;32m????????\033[0m\033[0;30m%%SS?%%S%%\033[0m\033[0;32m???????????\033[0m\033[0;30m%%\033[0m\033[0;37m.\033[0m\033[0;30m%%?%%?\033[0m\033[0;37m+:,.,;+;,.,+\033[0m\033[0;30m?\033[0m\033[0;37m,............\033[0m");
    $display("\033[0;37m.................................,;*\033[0m\033[0;30m?%%?\033[0m\033[0;32m???????????\033[0m\033[0;30m%%\033[0m\033[0;32m?\033[0m\033[0;30m%%S%%\033[0m\033[0;32m????????\033[0m\033[0;30m?%%%%%%%%%%S\033[0m\033[0;37m.+:....+.....+..*\033[0m\033[0;30m*\033[0m\033[0;37m............\033[0m");
    $display("\033[0;37m..............................,;\033[0m\033[0;32m*\033[0m\033[0;30m%%%%?\033[0m\033[0;32m???????????????\033[0m\033[0;30mSS\033[0m\033[0;32m???????\033[0m\033[0;30m%%%%?\033[0m\033[0;32m*\033[0m\033[0;37m*+++++\033[0m\033[0;30mS\033[0m\033[0;37m,....:.......:..\033[0m\033[0;30mS\033[0m\033[0;37m:...........\033[0m");
    $display("\033[0;37m...........................:+\033[0m\033[0;30m?%%%%\033[0m\033[0;32m??????????????????\033[0m\033[0;30m%%S\033[0m\033[0;32m????\033[0m\033[0;30m%%%%%%?\033[0m\033[0;37m+;::,.....\033[0m\033[0;30mS\033[0m\033[0;37m;....*....;\033[0m\033[0;30m?\033[0m\033[0;37m.\033[0m\033[0;30m?\033[0m\033[0;37m,+.+...........\033[0m");
    $display("\033[0;37m.......................,:+\033[0m\033[0;30m?%%%%\033[0m\033[0;32m?????????????????????\033[0m\033[0;30mSS%%%%%%%%\033[0m\033[0;32m*\033[0m\033[0;37m;,,\033[0m\033[0;30m?\033[0m\033[0;37m....*.....\033[0m\033[0;30mS\033[0m\033[0;37m:,..\033[0m\033[0;30m?\033[0m\033[0;37m....;\033[0m\033[0;30m?\033[0m\033[0;37m..\033[0m\033[0;30m%%%%%%\033[0m\033[0;37m;...........\033[0m");
    $display("\033[0;37m....................,:+\033[0m\033[0;30m?%%%%\033[0m\033[0;32m???????????????????????\033[0m\033[0;30m%%%%S\033[0m\033[0;37m;:,,..:.......+..;.\033[0m\033[0;30m#SS%%?S\033[0m\033[0;37m.....\033[0m\033[0;30mS%%SS\033[0m\033[0;37m.*............\033[0m");
    $display("\033[0;37m..................,+\033[0m\033[0;30m?%%?\033[0m\033[0;32m??????????????????????????\033[0m\033[0;30m%%S?%%\033[0m\033[0;37m;...,....+\033[0m\033[0;30m%%\033[0m\033[0;37m..\033[0m\033[0;30m%%\033[0m\033[0;37m.+..\033[0m\033[0;30m%%\033[0m\033[0;32m*?\033[0m\033[0;30mSSSSSS%%SS\033[0m\033[0;37m....\033[0m\033[0;30m?\033[0m\033[0;37m,...........\033[0m");
    $display("\033[0;37m................:*\033[0m\033[0;30m??\033[0m\033[0;32m????????????????????????\033[0m\033[0;30m#?\033[0m\033[0;32m????\033[0m\033[0;30m#%%\033[0m\033[0;32m?\033[0m\033[0;30mS%%\033[0m\033[0;37m*:\033[0m\033[0;30m?\033[0m\033[0;37m...\033[0m\033[0;35m*\033[0m\033[0;37m,\033[0m\033[0;30m?\033[0m\033[0;37m...\033[0m\033[0;30mSS?%%\033[0m\033[0;37m..\033[0m\033[0;30m%%?\033[0m\033[0;32m?????\033[0m\033[0;30m%%SS#S%%\033[0m\033[0;32m?\033[0m\033[0;30m%%\033[0m\033[0;33m*\033[0m\033[0;37m...........\033[0m");
    $display("\033[0;37m..............,*\033[0m\033[0;30m%%\033[0m\033[0;32m???????????????????????????\033[0m\033[0;37m..\033[0m\033[0;30m%%\033[0m\033[0;32m????\033[0m\033[0;30m#S\033[0m\033[0;32m??\033[0m\033[0;30m%%S#\033[0m\033[0;37m...\033[0m\033[0;30mSS\033[0m\033[0;37m.\033[0m\033[0;30m#SS%%\033[0m\033[0;32m????\033[0m\033[0;30m%%\033[0m\033[0;37m...\033[0m\033[0;30mSSSSS%%?\033[0m\033[0;32m?????\033[0m\033[0;30m%%\033[0m\033[0;37m,..........\033[0m");
    $display("\033[0;37m.............+\033[0m\033[0;30m%%?\033[0m\033[0;32m?????????????????????????????\033[0m\033[0;30mS\033[0m\033[0;37m.\033[0m\033[0;30m#%%%%\033[0m\033[0;32m??\033[0m\033[0;30m%%SSSSSS%%SSS%%%%\033[0m\033[0;32m?????????\033[0m\033[0;30m%%\033[0m\033[0;37m..\033[0m\033[0;30mS%%\033[0m\033[0;32m?????????\033[0m\033[0;30m%%\033[0m\033[0;37m,..........\033[0m");
    $display("\033[0;37m............*\033[0m\033[0;30mS\033[0m\033[0;32m??????\033[0m\033[0;30m%%%%%%\033[0m\033[0;32m????\033[0m\033[0;30m%%%%%%%%%%%%%%%%%%%%%%%%?\033[0m\033[0;32m???????\033[0m\033[0;30m?%%SSSSSSS##S%%%%?\033[0m\033[0;32m??????????????\033[0m\033[0;30mS%%\033[0m\033[0;32m???????\033[0m\033[0;30m?%%%%\033[0m\033[0;37m+...........\033[0m");
    $display("\033[0;37m...........:\033[0m\033[0;30mS\033[0m\033[0;32m??????\033[0m\033[0;30m%%%%\033[0m\033[0;32m???\033[0m\033[0;30m%%%%%%%%\033[0m\033[0;31m%%%%%%%%%%%%\033[0m\033[0;30m%%%%%%%%SSSS%%%%%%?\033[0m\033[0;32m????????????????????????????????????\033[0m\033[0;30m?%%%%SS\033[0m\033[0;37m+............\033[0m");
    $display("\033[0;37m...........*\033[0m\033[0;30m%%\033[0m\033[0;32m?????\033[0m\033[0;30m%%?\033[0m\033[0;32m??\033[0m\033[0;30m%%S%%\033[0m\033[0;31m?????????????????%%\033[0m\033[0;30m%%%%SSSSSSSS%%%%%%?\033[0m\033[0;32m???????????????????\033[0m\033[0;30m?%%%%%%%%%%\033[0m\033[0;31m%%%%??%%\033[0m\033[0;30m?\033[0m\033[0;37m............\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;32m?\033[0m\033[0;30m%%\033[0m\033[0;32m????\033[0m\033[0;30m?%%\033[0m\033[0;32m??\033[0m\033[0;30m%%S\033[0m\033[0;31m??????\033[0m\033[0;30mSSSSS%%\033[0m\033[0;31m%%%%?????????????%%\033[0m\033[0;30m%%SSSSSSSSSSSSSSSSSSSSSSSS%%%%\033[0m\033[0;31m%%??????%%\033[0m\033[0;30m%%\033[0m\033[0;37m;............\033[0m");
    $display("\033[0;37m...........;\033[0m\033[0;30m%%\033[0m\033[0;32m????\033[0m\033[0;30m%%%%\033[0m\033[0;32m??\033[0m\033[0;37m.\033[0m\033[0;31m???????????%%%%\033[0m\033[0;30m%%%%SSSSSSS%%%%\033[0m\033[0;31m%%%%?????????????????%%%%%%%%%%?????????????%%\033[0m\033[0;30m%%\033[0m\033[0;37m*,.............\033[0m");
    $display("\033[0;37m............\033[0m\033[0;32m*\033[0m\033[0;30m%%\033[0m\033[0;32m???\033[0m\033[0;30m%%%%\033[0m\033[0;32m??\033[0m\033[0;37m.\033[0m\033[0;30m%%\033[0m\033[0;31m?????????????????????%%%%%%\033[0m\033[0;30m%%SSSSSSSSSS%%%%\033[0m\033[0;31m%%%%???????????????%%%%\033[0m\033[0;30m%%SS#\033[0m\033[0;37m+,...............\033[0m");
    $display("\033[0;37m............,\033[0m\033[0;30m%%?\033[0m\033[0;32m??\033[0m\033[0;30m?\033[0m\033[0;32m???\033[0m\033[0;30m?S%%\033[0m\033[0;31m%%%%%%%%%%%%%%%%%%%%%%%%%%????????????????%%%%\033[0m\033[0;30m%%%%%%SSSSSSSSSSSSSSSSSSSSSS%%\033[0m\033[0;31m%%%%\033[0m\033[0;33m*\033[0m\033[0;37m................\033[0m");
    $display("\033[0;37m............,\033[0m\033[0;30mSS?\033[0m\033[0;32m???????\033[0m\033[0;30m%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%\033[0m\033[0;31m%%%%%%????????????????????????????????????%%?\033[0m\033[0;37m,...............\033[0m");
    $display("\033[0;37m............\033[0m\033[0;30m?S\033[0m\033[0;32m?\033[0m\033[0;30m%%%%\033[0m\033[0;32m?????????????????????????\033[0m\033[0;30m?%%%%SSSSSSS%%%%%%%%%%%%\033[0m\033[0;31m%%%%%%%%?????????????????%%%%?\033[0m\033[0;37m;,................\033[0m");
    $display("\033[0;37m...........*\033[0m\033[0;30m#%%\033[0m\033[0;32m??\033[0m\033[0;30m%%%%?\033[0m\033[0;32m???????????????????????????????\033[0m\033[0;30m?%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%SS%%\033[0m\033[0;31m???*\033[0m\033[0;33m*\033[0m\033[0;37m+;,...................\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;34m?%%%%\033[0m\033[0;30m%%%%\033[0m\033[0;32m??\033[0m\033[0;30m%%%%?\033[0m\033[0;32m?????????????????????????????????????????????\033[0m\033[0;30m?%%%%?\033[0m\033[0;37m*;,,,,........................\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;34m?%%%%%%%%%%\033[0m\033[0;30m%%%%%%%%%%%%\033[0m\033[0;32m???????????????????????????????????????\033[0m\033[0;30m%%%%%%?\033[0m\033[0;32m*\033[0m\033[0;37m+:...............................\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;34m?%%%%%%%%%%%%%%%%\033[0m\033[0;30m%%%%SS%%%%\033[0m\033[0;32m??????????????????????????????\033[0m\033[0;30m?%%%%%%S%%\033[0m\033[0;36m*\033[0m\033[0;37m;,...................................\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;34m?%%%%%%%%%%%%%%%%%%%%%%%%%%\033[0m\033[0;30mSSSSS%%%%%%%%%%%%???????????\033[0m\033[0;32m???\033[0m\033[0;30m???\033[0m\033[0;32m?????\033[0m\033[0;30m??%%%%\033[0m\033[0;34m%%?\033[0m\033[0;37m+:..................................\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;34m?%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%SS\033[0m\033[0;30mSSSSSSSSS%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%\033[0m\033[0;34m%%%%%%%%%%%%%%?\033[0m\033[0;37m+,...............................\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;34m?%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%\033[0m\033[0;36m*\033[0m\033[0;37m:.............................\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;34m?%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%\033[0m\033[0;37m;............................\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;34m?%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%\033[0m\033[0;30mS\033[0m\033[0;37m+...........................\033[0m");
    $display("\033[0;37m...........::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::...........................\033[0m");
    $display("\033[0;37m....................................................................................................\033[0m");
    $display("\033[0;37m....................................................................................................\033[0m");
    $display("\033[31m \033[5m     //   / /     //   ) )     //   ) )     //   ) )     //   ) )\033[0m");
    $display("\033[31m \033[5m    //____       //___/ /     //___/ /     //   / /     //___/ /\033[0m");
    $display("\033[31m \033[5m   / ____       / ___ (      / ___ (      //   / /     / ___ (\033[0m");
    $display("\033[31m \033[5m  //           //   | |     //   | |     //   / /     //   | |\033[0m");
    $display("\033[31m \033[5m //____/ /    //    | |    //    | |    ((___/ /     //    | |\033[0m");

    /*$display("        ----------------------------               ");
    $display("        --                        --       |\__||  ");
    $display("        --  OOPS!!                --      / X,X  | ");
    $display("        --                        --    /_____   | ");
    $display("        --  \033[0;31mSimulation FAIL!!\033[m   --   /^ ^ ^ \\  |");
    $display("        --                        --  |^ ^ ^ ^ |w| ");
    $display("        ----------------------------   \\m___m__|_|");
    $display("\n");*/
end endtask

/*task display_pass; begin
        $display("\n");
        $display("\n");
        $display("        ----------------------------               ");
        $display("        --                        --       |\__||  ");
        $display("        --  Congratulations !!    --      / O.O  | ");
        $display("        --                        --    /_____   | ");
        $display("        --  \033[0;32mSimulation PASS!!\033[m     --   /^ ^ ^ \\  |");
        $display("        --                        --  |^ ^ ^ ^ |w| ");
        $display("        ----------------------------   \\m___m__|_|");
        $display("\n");
end endtask*/

task display_pass; begin
    $display("\033[0;37m......................................................,\033[0m\033[0;30m?%%%%%%\033[0m\033[0;37m+,.......................................\033[0m");
    $display("\033[0;37m.................................................,,::+\033[0m\033[0;30mS\033[0m\033[0;33m*::;?\033[0m\033[0;30m?\033[0m\033[0;33m*\033[0m\033[0;37m*+:...................................\033[0m");
    $display("\033[0;37m.........................................,+:...;\033[0m\033[0;30m?\033[0m\033[0;31m?\033[0m\033[0;33m*\033[0m\033[0;31m?\033[0m\033[0;30mSS\033[0m\033[0;33m+,,,::;+*\033[0m\033[0;31m?\033[0m\033[0;30mS\033[0m\033[0;37m*..................................\033[0m");
    $display("\033[0;37m........................................+\033[0m\033[0;30m%%\033[0m\033[0;37m.;.,*\033[0m\033[0;30m%%\033[0m\033[0;33m;,,,,,,,,,:;;:::;\033[0m\033[0;30m?\033[0m\033[0;37m*,................................\033[0m");
    $display("\033[0;37m.......................................;\033[0m\033[0;30mS\033[0m\033[0;33m:*\033[0m\033[0;30m%%??\033[0m\033[0;33m+,,:,,,,,;*+::;;;;;:*\033[0m\033[0;30m%%\033[0m\033[0;37m*,..............................\033[0m");
    $display("\033[0;37m.......................................+\033[0m\033[0;30m?\033[0m\033[0;33m,,,:,,;\033[0m\033[0;31m?*\033[0m\033[0;30m?\033[0m\033[0;33m*+*\033[0m\033[0;30m%%SS\033[0m\033[0;37m.\033[0m\033[0;30mS\033[0m\033[0;33m+::::;;:;\033[0m\033[0;30m%%S\033[0m\033[0;37m:.............................\033[0m");
    $display("\033[0;37m.......................................:\033[0m\033[0;30mS\033[0m\033[0;33m:,,,:*\033[0m\033[0;30m?\033[0m\033[0;37m:,,;+;:,,:\033[0m\033[0;33m*\033[0m\033[0;30mS\033[0m\033[0;33m?+*\033[0m\033[0;30m?%%S%%\033[0m\033[0;33m;:\033[0m\033[0;31m?\033[0m\033[0;37m.:............................\033[0m");
    $display("\033[0;37m.......................................+.\033[0m\033[0;31m?\033[0m\033[0;33m;;+\033[0m\033[0;30m?\033[0m\033[0;37m*,,,,,,,,,,,,:\033[0m\033[0;33m+\033[0m\033[0;37m;;::;\033[0m\033[0;30mS\033[0m\033[0;37m.\033[0m\033[0;33m;:\033[0m\033[0;30m%%S\033[0m\033[0;37m,...........................\033[0m");
    $display("\033[0;37m.......................................\033[0m\033[0;30mS\033[0m\033[0;33m+:\033[0m\033[0;30mS?\033[0m\033[0;37m*\033[0m\033[0;33m*\033[0m\033[0;37m:,,,,,,,,,;\033[0m\033[0;30m%%\033[0m\033[0;37m;,,,,,,,\033[0m\033[0;30m%%\033[0m\033[0;37m.\033[0m\033[0;33m;:+\033[0m\033[0;37m.;...........................\033[0m");
    $display("\033[0;37m.......................................+\033[0m\033[0;30m%%%%?\033[0m\033[0;37m,:,,,,,,,,,,,,;\033[0m\033[0;30m%%\033[0m\033[0;33m+\033[0m\033[0;37m,,,,;\033[0m\033[0;30mS%%\033[0m\033[0;33m;:;;\033[0m\033[0;37m.+...........................\033[0m");
    $display("\033[0;37m........................................\033[0m\033[0;30mSS\033[0m\033[0;37m,,,,,,,,,,,,,,,.,:,,,,+\033[0m\033[0;30m%%?\033[0m\033[0;33m+::+\033[0m\033[0;37m.;...........................\033[0m");
    $display("\033[0;37m.......................................:.:,:.\033[0m\033[0;30mS\033[0m\033[0;37m,,,,\033[0m\033[0;31m*\033[0m\033[0;37m,,,;\033[0m\033[0;30m?%%?\033[0m\033[0;37m:,,,,,;\033[0m\033[0;31m?\033[0m\033[0;30m??\033[0m\033[0;33m*:\033[0m\033[0;31m?\033[0m\033[0;37m.,...........................\033[0m");
    $display("\033[0;37m.......................................\033[0m\033[0;30m%%?\033[0m\033[0;37m,,:.\033[0m\033[0;30m%%\033[0m\033[0;37m,,,\033[0m\033[0;30m%%\033[0m\033[0;37m+,,,:;\033[0m\033[0;33m*\033[0m\033[0;37m.\033[0m\033[0;30mS\033[0m\033[0;37m,,,,,;\033[0m\033[0;31m?\033[0m\033[0;30m?\033[0m\033[0;31m?\033[0m\033[0;30m?\033[0m\033[0;33m*\033[0m\033[0;37m.\033[0m\033[0;30m?\033[0m\033[0;37m............................\033[0m");
    $display("\033[0;37m.........,+\033[0m\033[0;33m*\033[0m\033[0;30m??%%\033[0m\033[0;37m:......................,.;,,,:,,:\033[0m\033[0;30mS\033[0m\033[0;37m*,,,,,,,,:,,,,,;\033[0m\033[0;33m**\033[0m\033[0;30m%%?\033[0m\033[0;37m..:............................\033[0m");
    $display("\033[0;37m........,\033[0m\033[0;30m?\033[0m\033[0;37m+:,,\033[0m\033[0;30m?%%\033[0m\033[0;37m......................:.:,,,,,:.\033[0m\033[0;30m%%\033[0m\033[0;37m.,,,,,,,,,,,,,,\033[0m\033[0;33m+*+\033[0m\033[0;37m+\033[0m\033[0;30mS\033[0m\033[0;37m.+.............................\033[0m");
    $display("\033[0;37m........\033[0m\033[0;33m*\033[0m\033[0;37m;,,,,\033[0m\033[0;30m?\033[0m\033[0;37m*......................:.:,,,,,,\033[0m\033[0;31m*\033[0m\033[0;37m.;,,,,,,,,,,,,,,:\033[0m\033[0;33m*\033[0m\033[0;37m,:.\033[0m\033[0;30mS\033[0m\033[0;37m..............................\033[0m");
    $display("\033[0;37m.......,\033[0m\033[0;30m?\033[0m\033[0;37m,,,,,\033[0m\033[0;30mS\033[0m\033[0;37m,......................:.;,,:,,,,::,,,,;\033[0m\033[0;30mS\033[0m\033[0;37m+,,,,,,,,,,,\033[0m\033[0;33m+\033[0m\033[0;37m.;.............................\033[0m");
    $display("\033[0;37m.......,\033[0m\033[0;30m%%\033[0m\033[0;37m,,,,;\033[0m\033[0;30m?\033[0m\033[0;37m.......................,.\033[0m\033[0;33m*\033[0m\033[0;37m,\033[0m\033[0;30mSS\033[0m\033[0;37m+;;::;;++*+\033[0m\033[0;34m*\033[0m\033[0;37m.\033[0m\033[0;30mS\033[0m\033[0;37m:,,,,,,,,,\033[0m\033[0;33m+\033[0m\033[0;37m.;.............................\033[0m");
    $display("\033[0;37m........\033[0m\033[0;30m?\033[0m\033[0;37m;,,,:\033[0m\033[0;30m%%\033[0m\033[0;37m,.......................\033[0m\033[0;30m?\033[0m\033[0;37m.,\033[0m\033[0;30m?%%\033[0m\033[0;37m++;::::::;+*\033[0m\033[0;30m?S\033[0m\033[0;37m:,,,,,,:;\033[0m\033[0;33m*\033[0m\033[0;37m.*..............................\033[0m");
    $display("\033[0;37m......,,;.;,,,;\033[0m\033[0;30m?\033[0m\033[0;37m;,.....................:.\033[0m\033[0;30m?\033[0m\033[0;37m,::+\033[0m\033[0;30m???????\033[0m\033[0;37m*;,,;,,,,,:\033[0m\033[0;30m%%#?\033[0m\033[0;34m*\033[0m\033[0;37m:...............................\033[0m");
    $display("\033[0;37m...;\033[0m\033[0;30m?????S%%?\033[0m\033[0;33m*\033[0m\033[0;37m;,,\033[0m\033[0;33m+\033[0m\033[0;30m%%\033[0m\033[0;37m*,....................+.*.,,,+\033[0m\033[0;30m%%S\033[0m\033[0;37m+,,,,,,,,,,,;\033[0m\033[0;30mSS\033[0m\033[0;37m:..................................\033[0m");
    $display("\033[0;37m..;.;,,,,,,:;\033[0m\033[0;30m?%%\033[0m\033[0;33m+\033[0m\033[0;37m,:\033[0m\033[0;30mS%%\033[0m\033[0;37m,....................*.\033[0m\033[0;31m?\033[0m\033[0;37m,,,:;+:,,,,,,,,,:\033[0m\033[0;30m?\033[0m\033[0;37m.\033[0m\033[0;30mS\033[0m\033[0;37m;,..................................\033[0m");
    $display("\033[0;37m..*\033[0m\033[0;30mS\033[0m\033[0;37m.,,,,,,,,,:.;,:\033[0m\033[0;30mS\033[0m\033[0;37m.\033[0m\033[0;30mS?\033[0m\033[0;37m+;:,............,,,+.\033[0m\033[0;30mS\033[0m\033[0;37m;,,,,,,,,,,,,:\033[0m\033[0;33m*\033[0m\033[0;30mS\033[0m\033[0;37m.\033[0m\033[0;33m*\033[0m\033[0;37m;\033[0m\033[0;33m+\033[0m\033[0;31m?\033[0m\033[0;30m%%\033[0m\033[0;37m+:,..............................\033[0m");
    $display("\033[0;37m..,\033[0m\033[0;30m?\033[0m\033[0;31m?\033[0m\033[0;37m+\033[0m\033[0;33m*\033[0m\033[0;31m?\033[0m\033[0;30m???\033[0m\033[0;33m*\033[0m\033[0;37m;::.\033[0m\033[0;33m*\033[0m\033[0;37m,,\033[0m\033[0;33m+\033[0m\033[0;37m.\033[0m\033[0;30m#\033[0m\033[0;34m?\033[0m\033[0;30m%%SS%%%%??\033[0m\033[0;34m*\033[0m\033[0;37m***\033[0m\033[0;34m*???\033[0m\033[0;30m???%%\033[0m\033[0;34m?\033[0m\033[0;30m%%S\033[0m\033[0;37m.\033[0m\033[0;30m%%\033[0m\033[0;37m+:,,,,,,,,,:;\033[0m\033[0;30m??\033[0m\033[0;37m,,,;.\033[0m\033[0;30m%%S%%\033[0m\033[0;37m*;,...........................\033[0m");
    $display("\033[0;37m...\033[0m\033[0;30m?%%\033[0m\033[0;37m;::::;+\033[0m\033[0;33m*\033[0m\033[0;30m%%\033[0m\033[0;37m.\033[0m\033[0;30m%%\033[0m\033[0;37m,,,\033[0m\033[0;33m*\033[0m\033[0;30mS%%\033[0m\033[0;36m+\033[0m\033[0;37m++++\033[0m\033[0;36m+********+++\033[0m\033[0;37m+++++\033[0m\033[0;30m%%\033[0m\033[0;31m?\033[0m\033[0;37m:+\033[0m\033[0;30m%%S?\033[0m\033[0;33m*+\033[0m\033[0;37m;:,,:\033[0m\033[0;33m+\033[0m\033[0;30m%%\033[0m\033[0;31m?\033[0m\033[0;37m,,,,\033[0m\033[0;30m%%#\033[0m\033[0;36m?\033[0m\033[0;34m??%%\033[0m\033[0;30mS%%\033[0m\033[0;37m*:.........................\033[0m");
    $display("\033[0;37m..,.;.,,,,...,:\033[0m\033[0;30m%%\033[0m\033[0;33m*\033[0m\033[0;37m,:\033[0m\033[0;30mS\033[0m\033[0;37m;\033[0m\033[0;33m*\033[0m\033[0;34m?\033[0m\033[0;37m+++++++++++++++++++++\033[0m\033[0;30m%%\033[0m\033[0;31m?\033[0m\033[0;37m,,:\033[0m\033[0;31m?\033[0m\033[0;37m...\033[0m\033[0;30mS%%%%%%%%\033[0m\033[0;31m?\033[0m\033[0;37m;,,,,\033[0m\033[0;30m%%\033[0m\033[0;37m.\033[0m\033[0;34m???????%%\033[0m\033[0;30mS%%\033[0m\033[0;37m;.......................\033[0m");
    $display("\033[0;37m...*\033[0m\033[0;30m%%\033[0m\033[0;37m++*\033[0m\033[0;33m**\033[0m\033[0;37m++;:,*\033[0m\033[0;30mS\033[0m\033[0;37m,\033[0m\033[0;33m*\033[0m\033[0;37m.,\033[0m\033[0;33m+\033[0m\033[0;34m%%\033[0m\033[0;36m?*+\033[0m\033[0;37m++++++++++++++++++\033[0m\033[0;36m*\033[0m\033[0;37m.;,,,:;\033[0m\033[0;33m+++\033[0m\033[0;37m;:,,,,,;\033[0m\033[0;30mS#\033[0m\033[0;34m??????????%%\033[0m\033[0;30mS%%\033[0m\033[0;37m;.....................\033[0m");
    $display("\033[0;37m....\033[0m\033[0;30m?S\033[0m\033[0;37m;;;;+\033[0m\033[0;33m*\033[0m\033[0;30m?%%S\033[0m\033[0;37m.;,\033[0m\033[0;33m+\033[0m\033[0;30m%%\033[0m\033[0;37m,\033[0m\033[0;33m*\033[0m\033[0;34m%%???\033[0m\033[0;36m**+\033[0m\033[0;37m++++++++++++++++\033[0m\033[0;36m*\033[0m\033[0;30m#\033[0m\033[0;33m+\033[0m\033[0;37m,,,,,,,,,,,:\033[0m\033[0;33m+\033[0m\033[0;30m%%#\033[0m\033[0;34m%%?????????????%%\033[0m\033[0;30m#%%\033[0m\033[0;37m:...................\033[0m");
    $display("\033[0;37m....\033[0m\033[0;30mS\033[0m\033[0;33m*\033[0m\033[0;37m.......,+.\033[0m\033[0;33m+\033[0m\033[0;37m,\033[0m\033[0;30m%%\033[0m\033[0;37m;:\033[0m\033[0;30mS\033[0m\033[0;34m???????\033[0m\033[0;36m***++++\033[0m\033[0;37m+\033[0m\033[0;34m?\033[0m\033[0;36m*\033[0m\033[0;37m+++++++\033[0m\033[0;30mS\033[0m\033[0;33m*\033[0m\033[0;37m,,,,,,,;\033[0m\033[0;33m*\033[0m\033[0;31m*\033[0m\033[0;30m%%SS\033[0m\033[0;34m%%?????????????????%%\033[0m\033[0;30mS\033[0m\033[0;37m*,.................\033[0m");
    $display("\033[0;37m....:\033[0m\033[0;30m#S\033[0m\033[0;31m*\033[0m\033[0;37m+;;;+*\033[0m\033[0;30m%%%%\033[0m\033[0;37m;\033[0m\033[0;30m?\033[0m\033[0;37m;;\033[0m\033[0;30m%%\033[0m\033[0;34m???????????????%%\033[0m\033[0;37m.\033[0m\033[0;34m?\033[0m\033[0;37m++++++\033[0m\033[0;36m+\033[0m\033[0;37m.;,,,,,,\033[0m\033[0;33m*\033[0m\033[0;30m#\033[0m\033[0;34m%%%%???????????????????????\033[0m\033[0;30mS%%\033[0m\033[0;37m:................\033[0m");
    $display("\033[0;37m.....,*\033[0m\033[0;30mS#%%%%??????\033[0m\033[0;33m+*\033[0m\033[0;30m%%\033[0m\033[0;34m????????%%%%%%\033[0m\033[0;30m%%%%%%\033[0m\033[0;34m?\033[0m\033[0;37m*+.\033[0m\033[0;34m?\033[0m\033[0;37m++++++\033[0m\033[0;34m?\033[0m\033[0;30mS\033[0m\033[0;37m,,,,,,,\033[0m\033[0;30mS\033[0m\033[0;34m%%\033[0m\033[0;36m?\033[0m\033[0;34m????????????????????????\033[0m\033[0;36m?\033[0m\033[0;34m%%\033[0m\033[0;30mS\033[0m\033[0;37m+...............\033[0m");
    $display("\033[0;37m........,:;++*\033[0m\033[0;30m??\033[0m\033[0;33m*\033[0m\033[0;30m%%S%%%%%%%%%%%%%%%%?\033[0m\033[0;36m*\033[0m\033[0;37m+;:,,..,.\033[0m\033[0;36m*\033[0m\033[0;37m++++++\033[0m\033[0;30m%%?\033[0m\033[0;37m,,,,,,:.\033[0m\033[0;34m?????????????????????????????\033[0m\033[0;30mS*\033[0m\033[0;37m..............\033[0m");
    $display("\033[0;37m...................,,,,,............,.\033[0m\033[0;34m?\033[0m\033[0;37m++++++\033[0m\033[0;30m#\033[0m\033[0;33m+\033[0m\033[0;37m,,,,,,;.\033[0m\033[0;34m??????????%%\033[0m\033[0;30mS\033[0m\033[0;34m%%?????????????????\033[0m\033[0;30mS%%\033[0m\033[0;37m,............\033[0m");
    $display("\033[0;37m....................................,.\033[0m\033[0;34m?\033[0m\033[0;37m++++++.;,,,,,,\033[0m\033[0;33m*\033[0m\033[0;30m#\033[0m\033[0;34m???????????\033[0m\033[0;30mSS#S%%\033[0m\033[0;34m???????????????\033[0m\033[0;30mS%%\033[0m\033[0;37m,...........\033[0m");
    $display("\033[0;32m \033[5m    //   ) )     // | |     //   ) )     //   ) )\033[m");
    $display("\033[0;32m \033[5m   //___/ /     //__| |    ((           ((\033[m");
    $display("\033[0;32m \033[5m  / ____ /     / ___  |      \\           \\\033[m");
    $display("\033[0;32m \033[5m //           //    | |        ) )          ) )\033[m");
    $display("\033[0;32m \033[5m//           //     | | ((___ / /    ((___ / /\033[m");
    $display("        ----------------------------               ");
    $display("        --                        --               ");
    $display("        --  Congratulations !!    --               ");
    $display("        --                        --               ");
    $display("        --  \033[0;32mSimulation PASS!!\033[m          ");
    $display("        --                        --               ");
    $display("        ----------------------------               ");
end endtask



task FAIL_PATTERN_task; begin
    $display("\n");
    $display("\n");
    $display("        \033[0;34m------------");
    $display("        | ┏┓ ┏┓ ┏┓ |");
    $display("        | ┗┛ ┗┛ ┗┛ |");
    $display("        | ┏┓ ┏┓ ┏┓ |           \033[mI HATE ICLAB!                    ");
    $display("        \033[0;34m| ┗┛ ┗┛ ┗┛ |    \033[0;32m＼O/");
    $display("        \033[0;34m| ┏┓ ┏┓ ┏┓ |    \033[0;32m //");
    $display("        \033[0;34m| ┗┛ ┗┛ ┗┛ |    \033[0;32mノ)");
    $display("        \033[0;34m| ┏┓ ┏┓ ┏┓ |            															    							");
    $display("        \033[0;34m| ┗┛ ┗┛ ┗┛ |            															    							");
    $display("        \033[0;34m| ┏┓ ┏┓ ┏┓ |            															    							");
    $display("        \033[0;34m| ┗┛ ┗┛ ┗┛ |            															    							");
    $display("        \033[0;34m| ┏┓ ┏┓ ┏┓ |            															    							");
    $display("        \033[0;34m| ┗┛ ┗┛ ┗┛ |            															    							");
    $display("        \033[0;34m| ┏┓ ┏┓ ┏┓ |            															    							");
    $display("        \033[0;34m| ┗┛ ┗┛ ┗┛ |            															    							");
    $display("        \033[0;34m| ┏┓ ┏┓ ┏┓ |                              \033[31m \033[5m  i:..::::::i.      :::::         ::::    .:::.        ");
    $display("        \033[0;34m| ┗┛ ┗┛ ┗┛ |                              \033[31m \033[5m  BBBBBBBBBBBi     iBBBBBL       .BBBB    7BBB7        ");
    $display("        \033[0;34m| ┏┓ ┏┓ ┏┓ |                              \033[31m \033[5m  BBBB.::::ir.     BBB:BBB.      .BBBv    iBBB:        ");
    $display("        \033[0;34m| ┗┛ ┗┛ ┗┛ |                              \033[31m \033[5m  BBBQ            :BBY iBB7       BBB7    :BBB:        ");
    $display("        \033[0;34m| ┏┓ ┏┓ ┏┓ |                              \033[31m \033[5m  BBBB            BBB. .BBB.      BBB7    :BBB:        ");
    $display("        \033[0;34m| ┗┛ ┗┛ ┗┛ |                              \033[31m \033[5m  BBBB:r7vvj:    :BBB   gBBs      BBB7    :BBB:  		 ");
    $display("        \033[0;34m| ┏┓ ┏┓ ┏┓ |                              \033[31m \033[5m  BBBBBBBBBB7    BBB:   .BBB.     BBB7    :BBB:   		 ");
    $display("        \033[0;34m| ┗┛ ┗┛ ┗┛ |                              \033[31m \033[5m  BBBB    ..    iBBBBBBBBBBBP     BBB7    :BBB: 		 ");
    $display("        \033[0;34m| ┏┓ ┏┓ ┏┓ |                              \033[31m \033[5m  BBBB          BBBBi7vviQBBB.    BBB7    :BBB.   		 ");
    $display("        \033[0;34m| ┗┛ ┗┛ ┗┛ |                              \033[31m \033[5m  BBBB         rBBB.      BBBQ   .BBBv    iBBB2ir777L7  ");
    $display("        \033[0;34m| ┏┓ ┏┓ ┏┓ |                              \033[31m \033[5m .BBBB        :BBBB       BBBB7  .BBBB    7BBBBBBBBBBB  ");
    $display("        \033[0;34m| ┗┛ ┗┛ ┗┛ |                              \033[31m \033[5m  . ..        ....         ...:   ....    ..   .......  ");
    $display("        \033[0;34m| ┏┓ ┏┓ ┏┓ |            															    							");
    $display("        \033[0;34m| ┗┛ ┗┛ ┗┛ |            															    							");
    $display("\033[m---------------------------------------------------------------------------------------------------------------------------");
end endtask

endmodule

`ifdef RTL
    `define CYCLE_TIME 20.0
`endif
`ifdef GATE
    `define CYCLE_TIME 20.0
`endif

module PATTERN #(parameter IP_BIT = 8)(
    //Output Port
    IN_code,
    //Input Port
	OUT_code
);
// ========================================
// Input & Output
// ========================================
output reg [IP_BIT+4-1:0] IN_code;

input [IP_BIT-1:0] OUT_code;


`protected
PCE?I@=N1L@YJTP;VS)DD),NdNU#84SQ8AP>aV+XMDOX/^E3P]GZ5)UN:6AO=QBS
a90]db^QgNO\_N6>F-Y4J]EF3ZH:P#(Ne_/+2D/5GI[W2YO=D7J1f:gH9e5J=1M_
L->6a#MQZ&8QdQ0B2(VA1<FR\9H3/PQ10<L,bCNGZX[0Wa>#5Pe^dKK#(NB)[Z7J
?d[=aa3G2;c8@42GQ;:A-\geGEg8G/?Yf>Y=D;=;3gRFIgTT6fffV63/4SdVR#>S
0&b5^GgC05=@5M]:9RG6D(TbLI165@;A4MM+(gWgfFV8L:1^(5V]:Y>Z#7FBB/:.
+T?2gYg@P<#^+8cGMDV_,.R.Gcgc6Z]>#PJ2ZQJMOdb:d>RD#+Q5;TdMLLE\/cH-
(F^P/dLRTLF(e/R5_/&L0#:;#NL0L)fCU[T-2b^S436gP\(6H-6R,YTB\BO+1SA&
CEQ0=LOb\@=T^?MV,B(#BMY?=5]3Ib0BY(<=\ZPVY]c;0c]7CV=WPC.:GD@d0&.,
XV,4.2_3BH&]@]M6?P.-9aaH2PIMf?.7c8,U\)a-RAUT,JF^VPC?1Z-d<MKBCfF&
AD4DcH^@A[WJfgP\DY1-:Z7NBS&89\W-TfH-b3^/7G9>#AbaT\2BH74SH[W=QG::
NNRbeF_cf+M4@6G(YBLFI1c4X3&HY9#fL>3M3Acf2KF79=42-<(3fI9M08L9+0cX
C]ab06>0ACQc=]-MX&gAH^=#OD5Ff8H8R.QF_6/T/N4W2#GP3XSdH@2^]73^;N\Y
_KKRK5MLG^/cK^)b_?_WaM]&)<g,5=:N4D92]YG>)JXCT0ETQ_If^.<1]X>/5eYM
D^0IP5QLNABLgg#:.D\gBA&P/5#YNLM_c[\ag=QNG^-I5Se6Va4d-L#/DcY4bg/(
KL0TfH)]U13cQYQFS>A4EKB3HM+Le;P-(BF8@XUY.>8ZHJ?X+/+?^8Q\b_<MCJ&d
H,1=EL:&[4,[(CKR:H(@)UGS8R8YU3[N7fX@7Z1K7G5(S]K38f/aYb8/>URE&HI0
R)<6]01-A9e1aDN\EgPV)@#745e]YUV&g@3bYe)M<UaOZE]_X9=EQ-c?-e[c[983
1DTE;/ZV57+._b0:.M^L^07@9UKGC<.4:KPX3]O9P[+DG:501KW+aHV)\7MWR9S0
X\MFH/C+Cd@I5=I&]?JU<J]Q-eTOgeEFNHP4DV@2,IWN,EC&E:VgXU3SU]]1F6Q3
B0BZ=TfG3=XX_#N<>+CYA#M\0=E&a-a>ZKDY(8c4R\L6P:dCA8K9EN3L?M^:T_,(
PSC#HU#?<)8BIFIDTJXNNA3=\)X/\<KA\2?EEf_H7VM<?fZ_V_XZ[<T-]<=9?fGO
Ha6L2KYW0fK<YQ[&PSSb,L>BJOW+Pb1fMSOEAdbEfeWH#N;P@I&56>N]#d7=?2/9
R79JS&D5ZJ>;aTJ]9HEJ\CJMK).Ef/]&2a:F[3^6H)CS&K5c#(F./8[0)U2ED(#,
N-b/daE#gEZbaXg_6eLZ@(:7f.S())WL82IVZDc;L<#FMgU+-c.=<_3T5]TRgRF-
ETT.Ba=T/5@G4XG-d.6:RV(5O7L.=]N3+Ac?79QJ9A3U/f4KA;^H751EQG.MJU;/
F,e[7]#W8+S)=/)G60F1C-2V@aWRAZ#d,/VOF:]@)YN[:]@>36Pb0ddPFSQMBX;/
98&Q>Y)P<?.J1:5/.]\0\GcVX?@E#2)3-JSgT6S;TZLHDLQ#@PCaO=.P8Ld^,)[5
]g_BHeMIA5UY401?,Abc8/J7HSF59cff@,AV)@OD#=K7bA0S5d[5PFW_LGE6J>#b
Xg;CRM8Q^+M?O;9S^?#YbITg6N29;^GZH,_TgGeSJ;=?:a+MHZfK\Ce4\A4EWfEB
W/b=-I0aecA@gc(AbZ:XXcX\^-0g&)/:I5_P4QF9XU0gHW=CBOe6^.(eC@NIF-IY
V4dO2e-:IK/LV1Z>UOcV=B&F(.JS]RH3eBE-;d5bYHcHARS-83g[\SQ>c50d0)38
MNQV:f>&>W#(=M@JEC_LHX\+^1@(61?]Ga@;Y_=[LV;\>L9.2[4H.H>g+E9//8MR
8LYfC5RP-6\D?+9Nf/YJ709Y]D8bIf.?NPf^X<D:f3#^3I<R;ZHUQ7(=V6CQ0V5O
G>]29XZXZP-V5Ac8S>g8:D\YA@a0g5AQSVIH>NVB(g&bQ^AKbUAc80eM]aPS6Z7>
#\I;AR?>2:^4K6G1][.SNJXXR@PM5fFCg_3<4;a_@QM_H]ed/#)DD)2/:L0O\(1H
OK[(S<0(^LF<gI7P8Ee@e)>YOI(Q+]B77Q;H2gD]^/^a.fAHFeEfE)/_(G\]7@4J
7@EOV+fL1WdJgVEO_[&GKb_g96KdAXI,9N]5-.&1CY]4_.:<W8LPT\&7]QKaANS5
R1<&F@\:2#AAWZ-:>>Z(5g@O;?<;7_dG0DVJ<]4Dg^[-.DPK1>fd0SIF6&]BgGOO
&.UIJNNGQO+6c91eO.d@36+^SB@W2XW&LI0^TOa;[14/5=I^9D^DEI;X76_TNAM9
NED#Db<>?W;;1DIga8N<F.B@0gMC8MFZ9HMB/a#P1..M?f(8#W:5)&-^VKFQ8g6;
>:5Y#2I]X=be/V4MA57CR=VO\<FJ2Af[<Kf[.5^P</,#L?J/]VLg9#+-b3\OPMFd
C;WM-V&c37MT+@EF4dD_]_?7RNgE6N6&Z9+TZAXf:1.@GN[EQY_4SMBA@D2LE_?Y
dNLg&-3V/b-HVC:F-P_XRKH.+Kga@[3[XZ-#7#&9,K#MDE#R@<TK&9@WH#SbS53G
&-YN^e:f<,7G?K;212>H#4=?7>_[:ZIWA(\FgL?2Ha1TK/f:PA4T<H?.,6<,6C?g
HGAX=?-XN6e5J[ZJfNZ<-(T&6R<Q_^Ma#4,F&R9aTNNf,B)E8U/RF-1FW;D3Ua6H
XGY,[;gbL-52>?ZH+.ecK.V:@?I?+g<cPZ8<46(\X-;T5ZR7(KQ61JYPDTF?ZeIa
3@<>Re,N#L0YbGR+ARN/+J4KfS:X)XQZAMe3H=;;Hg]_@2Od8e5PG.TW9WQa@-W1
_K4=@dYQD8J<#NTaT/C1,E0O]>4)UN\Y,R9<L+R9TA3&aHVAS#gHH5Z+X[WYSRQ<
^ZfR9(3=(GNgdOUdRAEYc?0VP3CON9SHYG@BJJM.Id7;d[bA0LT6S_b_([&@ce:C
6NS9a[9X\c5d.A\:8&UAN[(P])L-e?:XFMb?fSV2O8HI^.f9V)(FH8@?EATO#:FB
(B\JYA2W?LSR4>6K61RQU_[FM:^=]WJ9e2?6Ge<YQ<<aNSf_#9M\=Y8@\aP7^eK1
^D)BV4).OW9H5aK^4^K2IGQf)FRFN#_HL@]LSGK<9+4C(b.e0e9V5\OEL2>7&V0E
a7CEdN9c8#IIdR3QH,OUaSEeN\NWRc/;@\/AeO:VcL:7>cG7)(I?)g73e3S5\OEN
OTSS.O:#KKbK1eH9Q/;E2XaE02[-P6e8-GVU6cbY8_Ub30b\\]gJ=RPNbOg0P7#e
C:9WagOORMZL;]a7J,&AdC#PRgd2X00\]]+]E3c_^4La@F>DWVa03EGHQDIH,U>+
/W:/H(#]=N;CY;K:NG&JB)_]-DeSIf.4V<U=IR;T[-Hg>G]I>D-MA)Fb\d>SOM[@
VP]>]_2+a4)E[AWD^<?\T,b;)A;VIaEg]BB()JL#[RVYab@3]YBZK0?;J;c<AXN:
ZY_XJ#+T@@.N[Q<_PE070&+)XT&<d=X.I73E92Pa_B:<?B2(SU03MZ)e@OfM3HUK
?;HaDUHWbceGSXAKT(-\g\D4bg&T+E3.[(2YG9?3JL12U\._[S9A><UM/N9911cC
CV_KS5&5)D^a+7Zc/29CU5)CK4TKL&^6+-g&gd#IH3[=g+ZK>B#>?#6Q8;b\^0V2
3^f^([W-Z@dCUE_@PKH.0fMO+eF7/c:N?^L4._6B:MCT@OB\gD^.ad#C^EZTb]Of
Y7\e/,4PEQ/6D=LK_JF5XUSRTG&0T:&;YP&.Q[0<D7M<Y>Na5G+13N]ZF2O;DD>c
(DB;d)LOL9L?5McR[Mb.9IHIE4<YL,]81b@6UO+9J]-&\:,H=e?&=^41ENXT2a)Y
+2HD?92fL2SUc,gV)bcM;]#:4HO-aT4(4\D?M/&Y;>A579\g0E-[ZEb5,9DceaSM
b#4+,:6<Y,7SBgW73@T0d<&)X:gFA#gKE<QYcC?X08++RCb-KIHS+4SV.RA.4,[f
3&+@4V?K0f?MED5UN9Tf22#W]H@/CNN8f)#2RgXQ=,#X=3.A1(5Lc\O#ecGN/.ZP
0B<d0RBN5V^TYMM#O?WXH]:NB#EFR=HYI.AR;#73<N9A]V0f4ACJ2826LROH3[VX
C4eI?_CJ?5)aNTLY+<FSCAX8^+#(If_6@e-AHYW[I\Y\JI08HI?4#TB6c&5X052H
C[R3XgN)BC^&-/73Q^8L+6::__0F?]TT5Ub,e-=]B;R+3E.HG47ZH/CL@9cU/R^0
J-dATH[-64SeDFe]5WC8>.Nd()c6?Oc1NdQ&?Xa3f)[C.)+/\V2/d[F(5JV8@UHO
LfK3\&K4;X:c.WGPC(.,Q+>S[fSVE3@4g6]^TPRD9MS/)a&N?^9g&3)WPY\=>]HU
U@a7AGgB+.QYbL85,&OO/5TM7dW>UG1#2IM4G,4LAb2+W[F9H:DW,<3>IA9aED#.
XS8?)(&d],DFN?GA#-<-5N-D+,MC7BB7XB0)E/U#RcW7@dU(3W49Gd_K&&+?X(@0
-,5?.e)AJWVD4Kacd3[HH9RD3A;D[>R+LA0e6Y)N\PV0d&X\cSdD@RLb1Z6#2QQ-
G/11:DR9g<,;[SIcW=c:>/?63Q_-bHc6@[/@P9GO,[f&1g&fg[ZgGOOFHILQPcDH
(+)T#9<T/RQeDVgJ70gYEO++W(&3)?NgFg=D#=_3aGYH<QP2=27SW[@7)+-Cc.\@
cR2.&a8-+YgIGOgFAT16V9?DCA>W@CQX4]EaeMZ:U-dA;WX(\A)e?T\2V5>Nc16:
Ya5Hf@XVP(_Ad-Sb/??(XVaKeRd_UP^/@)2g1\f9IA2fcHT2;&6ScTaVEF6f[_N-
BN(<b##=Y>/5^6b?3P@+U<eD,b5DC_4OI?VVHQ^SM+@CQP+K#1D@FRI+]<)(6dX1
HI5U)A4b>5L?NBOLA_gULZLaGA?M9[fL\E91<<D4fE4I>LA)<_G(O>OS7T11U6KD
eFG=ELa_B5Ae1L#IU:J,7c_QAgId?gZ2gFQa>.Y=J#L4d&+;25+Y#[9P+;OG2]AX
Ie/J^DJY9=K53G7]RALGJ2+0\9#RR_U+V3_CH0eK8(O>g#9.SA2d#Qf00Ie]Og34
5M>a&8M_=#HX7UcQ.NUBK6_5U3XY\KE;^]:T88Z<_-^#J);IM[B32,T6/5GEg8Q)
Fe[H51<TT&0QF(-29Jb1N:K=0[[.59/=YV@059Yb9)QK4B8[SEa=QO-L-QB5)2^:
&6KU&:QQ(^O9B-BaJ^g7>b?4?KP,V1@212YgMPX)PRQ)::N/9J.fY.B6[U.>5AgX
)K5\Md\?cQ<@2K.,_=U3;.JTVK#bV-G7]P2d+;F5A4eVWQE=2OB1-B>DXNG480&c
TG]cQ-7eLBggg1IG(RLQN4IM8<JC1\/,3:gT5_)N2X^,=7EDG9S#2>362MIL1LXN
T)=^+VB=IO-W)V,<F/#-)>_M7TR4J7&>4<_&7bR[0WD?==0d50?C^_-&-<)MF?70
&FZ[]1SF9F:__FZX?UU.ADDLV]XORBdJO24QQW23]d?;N/9^L;[6a&8>)6K?f@17
-,I#TWD1_W;OPfG^K9e6;U#/d:?H&>IWSYE&d9KAQeI7Z@3&[CV[g.&1CS#QDUJO
XO:R7DLG=I-[&G+a^EPUOCYD^6BQ(C9/&U_9^]PB71IK>.V@VMATf0\Jba&9Kb=R
E;8^Z0D^6^Le.G9U?43<@&2B:N-QPfS0=.eG\0KWf;PCaLgNb.@R1;2AB+-C&5AM
R79YSJW1ZVG_fcU[Re5.N^Q-Ta.Y^V_D#fTFd#85/8AI_UD2++[dF<2fC493YJ^#
0a)\?1F[7U9F(3V^\D:,UI[4f]3fP?U6(gCXZdQ47WC:Zd2_,9EV8g/#^[0f-Fd\
Z,[fIBJ\&)\4T.>CITf[6EDMH_b@/V;8Y0NNSQYe2X[bb=aHFM8TNfK)A>BgO_cb
)EXDd/R\&FQgT,&IZfK3-b50>BEI6/Xb1Ld&8GL2^BGe]aQfHaJ:&?aK^CM4[FAD
S?e@G.5PFP/7e_\^>+#V@S(/TPUBKaJddVLR=36<CZ)B81cX#EVL@AAF2Q2GaC_I
RT81EY]WQQe=,QL,DW@D-&2=3SBKb^^-c.JQ?S9.CUGaeM6Cg]W[IH^2.Y[b)7Lb
H3&L3aU<</.]4HCW8(g-g&C3=(XR)c2/RV?0E?IR9Vc#8VNf=]8A)S\310&5:VTC
&bAbc8Qc74QZ].LULZCBN0^Q2P]\[/9.Lf2HS_T@efe7;&+H;cG_B^d2K]]H6b/6
Fb#VPF8,\cTX5HS&4f7P/db<OfI&Ad35&QZRgdb=X745E4\b?4K4+aTJ7DN)4.P7
E-0ZCX3/,5fH;cf7#eMU,=fYZU):Ra9DK.cJ4fP&>eN<-d;dTE5Ada3L[M=@W4Y?
)@=Vf=/RVGH[GDA&[8F>(-Y,,P^>XONAX>0Nac_DgT:b3AQ08g\g&)WS,:PB70\O
U-487@BbC@=CXAW85JOG\FW>J9/2CT6H^R;_H&7aJ+Q75E@ENB-\Y8?a?S12_4HR
ObDZ6Y&>D7X&G:]70CS8c0BV3\[PfM),c.a,;J5L\#OMc[B34&L14>8]P^VB8I&Z
bV1AD-\).K\>51R=Yb&(Ha:[[fc]WBf79)#:J5IG8Q5S?UGLO0CcHRf]62A,P4Nc
^F<KKc52b11@+1A:VV=CT&TbA8H.GHGPeSJ;d>9EX0g.:U^X/I,>#Mf\.f?2VQRd
Z1)[;SaPJCFY?(#;8PBNZT]=DZg-UaSC[.U/-XW43Le?eK,Q7E&Q3&>_]BH=ZX^_
[VFHY=)JHf/9B-^eSCW#/AVRU2e57J6&[U1gc=/dY@^#,5)75+#3\B)DS:E<4b_O
,?HKWB18<b<QaKS(AB6DXfE#ZJbNg/NM4U=bL=T64Q8,.9AI&&,RMEG)K0F.NG:\
94YL#eBU7O>H?_]<O9Q,O/Rg@>NNMN#78^XaRN1ET0RC4KHBa8Wg&AJ8VPFe\\JK
/HTSWQ-cbbNM@<#6g-D1/_PD<7K5XZUTE1TWd4TdA-@CR1\,WVC7bK=VUAefE>7D
4Je5TLHRd8aML6ZI\/2/U(13#+L74:C26D8)+(D@ION59.JJ->LffgF39I4fZgN0
<CIFE5_Ag#(H^NE:gW5+KO+UOg0J9.I2/bbKR01[:PKI6-()F77B-d/f55+>O5YH
=eDKX.c<5fOR0GXOCQWSdLReA]KD\_[feAg?/67fg1+eS#P7dQ\#/SQ9CeX<-^<>
UEPd5U@GJ7FS3P(0^8g[a>bg/R<R1=T-c8CVAf9^H]9KCY+&I647NI-L1O0&M#dE
g+UcOM^_D39;L.9)f\<Yag-7YDQ[08T=c+dQZ>T>+/VGJH7XHAADHfV^7,UT8&2\
e:CG/,cX:6#(GSJK5TKC[<REaRL&-AMRT;-Ue4(cK/CJR;H[[#CY5BfC07_P([5a
O(.+#16;)YGS#U6PKR=f>.c\JaN6[Ge9PPFBBdbZI^<0U-E#3=JSOO(1ZNB9VcHT
d@L.I?FHZIbM9SF]147a0.f96NP,+EXNVI\]-]#>VWD9X>G=M[]U91Y.3(O<O6:U
(+:)#-#\0<7HBJ2C6/=Zc&OQ7.]U-]M@:b,.I+7eOHYS3AQW9KT4]=T[8WD6ZM.1
2CCZO]EGYf2?=J>PDV0,5(>L4UM):1DWKdV[1gL4)(WHWLG[4a]N_Y5KT:H,9\NR
2G^cD>GF?Q<.AVGQ>1d[_#>K]:YJS)b<MYRJM,F4/]SY]E_[IJdJV/&/Nd//2>.]
QLFIa)7O0dAHHZQ<0+M\eRM7Y1UF(=C,PJQ^ESgVIOc=-N@N1X].H@UbL<d8L4R9
GL]9IR=_7:K6/_(+GKFC(;OKb4_+D#+0eR>:H8=BXHDWLMI2^6bW@EQ=d>NE(:(?
6BSRN[SKFY56>f[WP9eDCOCTWUJ=;CHYGE3<RA(ZU_8fBEF\c#IY?NED6[ETOI-<
:?-+EQe;,P:9OA9=B.Q(eS8R>FDbY)&d1=5aA2KR4&1H.&H#D,N=2a0GcA)Fc_M[
@Q7MZN4;0/TFdAb?80_b1.E^<F2Ge;KaW2#<G[Y-JaOAId#Ze-ACKUD&.=aEeaG0
L:H;F:/-_/TO\#9E9YeN6Z#>MgbNeW<)QCbFQBaHF/NENG[g@8OF=+5aA9ZH<F;V
HJJVTf(WBS8SaVH8DfVd6L1b?IK?34C]TV^Y:Z0U)ZTCSXG1A1bR89,-NI5.W\KM
^J&&2Rd0Nb(\dCaM8LLC3>8^,E?9Y9@9.B.FY[@TF0@WJUX#C)J52<K#:Y<<#.8;
W&/Z)U)KWHWg.,3WeJVP;FSEX@HC.7)M(YWO4VaD>-cF:[JTGKOSa/Q&U[b<WJQ0
-=X]DX\&6-(_,2AZ?0GaP5f9^6@=&_K1e[R#VI^)31JU+2J>2ZbO[&fV<WL;W63I
Q]b-3W9d5@]J<VS>L@K3RTVKXUD]E(IO<>YYJ]E0(5QQP&\ULG06H<<5NYPB3e-8
<3^>H@HRB6^[85C5dX^8?/b4E1VGFN9RAQd#SELaBbXERU/;9/2;VJg4A1bHW,ET
1a64S+e(gYLa]8^(B]<0WgS2JgA2(?Y_Cc4GcOCU,6#(Z@L;?312/K>M+1>:=:d0
a2F^f]fUL.0]X7\^VAHf>^F,K^I\&7gP.aVK+9[-RcK,MRgEEUERaT=SEF[I;..R
d<5=ZWPZ4?R;MJ&CS<P]-N3W1GBX:477DJL:TT8A:=DHN;#TMDT-OI=MZI(Wd1@b
Q-#<M7Yf;@LLYED<7\b2:+-7617M_\WD45-S49]QU05K>/^]/4LGeQ&gFHZ]F@L0
ASP(YQHKK#Y1B1b6SaN<A1bSPB@3I9f[U11DeG)OOL>NMBRM&Qc,7cfU1Y-F?.-+
.KBB:0RJb1)JaU^I]+Kd#=.1+bH8M[G(FS&eBT/WNBU54[9)KK\B/5I]P6;0)JEd
+F05gV>832PCZdWO7>Y;17>_5a[e.-ASI&A)YZLgB;3#DegH6#G-+N_:8HJ[4H2g
O&?5fd]dSEA/@I_eg\OEPb2R8N8QH,aUA2f]d:fGM]W+eO@FdaB6==<Y9DGJM:Mb
5&/#fBHSI\UQ:_dgW+A4/Aa34Wd9&aL<DJ/f].9(M9aW5I3/[;<=[K:P,);YCDVf
]_gID6V;W;-<NBgY(CK>GMJ(=KII)OY&KS;RTDcbW/@N+1^U#1g&d=A+_TD3&(^H
?TXLP^W/Z?Pc_<-GQb&1NC;^dU&6DTA:/0J,/>K)4Y&42b[dQeX48O/Q?OZ[)-d0
6LH;[9;4&8);((:=1DBUEC]\PMTJH)IQ5cJTAN@JK[C4AVC1WQ7Eg+72+WeK=[b)
^&C<NB3W?Sd+K8XTGR?7gL9<)+A7?FYbP()LXI#Y5T7814SDA+J[/0&K3Lg\5JMG
Gd2-1eAaD11F=Pb\G)NV3V]Y75UO6<0a[AK?NBJK-gUa/QUf^(dDS6OM(#_Hg^[d
:fd&8b[2?KK_S.\g]a^@19@gUOb&0OBH+3NEg(G3-4(dae?aX4&\@09+Z2D6=OTF
=[8C]EE+S:_<d)LCO>JEa-W>8-9,EO2:Vd6=a,A?2)aR[-/UC=UaJ@+.#7NOI8P<
=Y#+VM&]Z)?/O)V&<=V.7[[P,<5P+QJ5H>AaTI7GY7f&,=6I^cFY2),fEYY0BX:I
(#[Z5N\DI+@HF?,\[[eP?9BgC@77]<-B/CHNad7?3XVOE>:d0#:W9L0>F-,/@P,-
Q3b,c3:AF+<K=XR5a7;K.6\^LFW8[Jg;Zg&O\)V:97H1@aSLL7?C>39a.cZ<(2YS
&fJd0.N=G)Ma;1MWF6.\J-QH)S4U6A][A[NX+_]0JJAKJV@W6544(AE(_Y@Vdf:Y
J2^K:.Tde&^,8A3]<_4UI[A:d.J^NL-cbaBR_Sb1dC5MNQd#C-X&]CA<+7Z9&(72
]6:1#;MN1)-UdZ0UXS5_1]:VQK989N+]02@72>RO<=[503=;&?:XO\g_@-e,R-E#
XOeG=\J>2=J16dM#Ngb5McX76?Mg]9RJR@Le+g;L?(J)99K,)KY&4aANF4c0:9Z@
CIP-\3^R9cEIN:Q(S8V)JPMFOW)e>N-Y;aE0_ROG=X5FcFL4\c,:L3GcB?.#:e,8
Mf0./756HIPS?5Ag9W]6b:P]UYcf8UAb-:P32Z>J99;8)YP[1.>_4cK#X;g5Lg_-
:KaT:6H:P>S[Wa+W2ZD6.AN)?<CbUP-KN@W-EX0/8RVPbUCP[)GUUVDGH;]P(K?0
/dc8Q@.,\-TOC8b#f4H.E=Qb>867VSM1f059EWYaP0H)a;3O52CA#6TZ.K7eS?72
W@2=Ib2)g)B?A_J4-GdG^08N>\SAUVHZM&DVV#SAE)4YG:K.6,ZW6O<G)93.D1Z8
1(W@V9YJ<7ZTK6Ad6_>eJTAVGO+\>/1XNBVMV4R],QaY@R@3g+Ac\6=[38g&9M;Q
f_BJKXG2L&P]A)T8eGE)56gMGHUZQC-G+C)_UN37XVZN#^LK4U_RP@7UBe:+cOa5
2DNDD0GZb=Z;Xgf>H=S8Q&(0NQ&6/?@3VD(AE_8D#T8UD?Na,Y3<85F7VZIYeE6X
ARX7R6XD-.^ddE3(R7\\_bVR72Z0&fVQ1+faQ;dg,EY/H.DFUR@A)R@LaQ:4fcYU
2U[+?:8Z/K07C&(HfQ,E^N4L-)62M2fVDYa+ERbEM]2(E+@]Sd]eWbfb<F85)(D]
/-JY2g9PC]NcgEO_I^UZ;S94>42WK87_N.4Z-PdaVg(:7(#.PVE=WD7<T:Y9>T?V
AHR74DMWF30B@,E48@0E4HF.A10MGDZR;3:DPO4#-7;XbU[+HE1F^74\&_Z[-VC?
e1cN(>R<EWaD3J/M(&O_JeODe[/&aQ(D.Gc_b#HEP;Q)>;VN[6gS8VHJN6gK:1[A
[;@EL25^Od<UfEGfe:=O(V>gLR5VCT2444_ZcYSW7@_::.?\>&\8J-))=Mf79&/S
,WAfJY(+S(a+L@.C9KFF4.O(+(.Xf.?9S)U_GM8RfL)b;YWVZ#2)GVM80aE[\A87
5-#/N3NYH<Y.VQ[;_d4)Pge3+7#?UeZeS11.QKRCF[S=J10g.QC&=9K#,CX)VC0J
9T:+7+eN[^dEc0\Pf:W;?9W6Rc(Y&NFJ3g/KXTP^FO;162@V_fPeI&R?>G?VB##[
(1bJ24-geK9V>RW#((_I/-O\2Ea3<V8:)b-JbWQ2_<#,#590\QT94R<ZC_ZNXK-P
:3#VbQX10/)TST&1af6Q^[_;?CbXD_:-(5GD);CY<252aO[AC2aNSWO-5L^3a?cb
3VQ],?7OHYW30J?Y3:7GUA9N35JBXeJ8?g<5[3&P(gYc]?cQWDUTV38-A4#5A7FF
+SNP_;]OaEIHJI.-M431^aNZc>C.5Y=[G87_L]_MY(@JfD3P)04GAX>Z@T0+F321
-8+U)A:D6/\KY[:0YeYW9X]BX[=25;5D61EL5CR<2IM=+FN,+&>FTN-]B+RRb4IF
7TaBQ]bBETZ>RR7BZU?J8]+GWYK>QM.378FP5[D23bRfRgVc5NfdGQKbaQW.NE[9
cZ(//ND;GHI2(X@@S-(I4G>QX/e/,\\A;.G,VadJMK@a.[fbNOB;6eT-1_?GF[=Z
)OJDYQ&>O]VXCVP;FVLMB<<KH7f@>O4IG:KGUIW]gfU:4CKg_QS9Z>1>?1=OUF+.
X9=11UF,]JTHW7a/.IA(QNVKfT0_>PN3N4+T3[e3K>@#2Zg[)&J_G<;_6C:YVEbb
7E6=4.;b[XGJWPWJ^V^73NC5^AG#cIWL;a=)4[C6NJ88TE])IB<O[FGRA64,_e1K
RAUd.S)_YXQFb.R8I/>W20g3^+H]HI:JaNPg@e(3)E0gLYB-EDQad29OM)\Jc&9,
O1BeI0YHZ95WT.MLZbGJWX^;)8N?TT_V:aL=MK6&\S^N]](NS:3BJJR<9FD10__(
#/3N=\74.#a0#V-O2)V_@2817:AFK^N>9=3WgfXB>#BFf[-H)>UX\5;SF7H._KGZ
@F@dTA<N=9+cee07T&-TO@E(E:=Q,M23b[SWN0OA2@f[KHF]A--a.=(N9.0IG6Hf
\#C9b0.0Q&KCX:?+XG@dgT>I87>@\ODQ8X4/d.)WY9PK^KSPB_<+J_/;)cVX7]09
PF^=9KWAZ:D[J9++WdV)+6(_64:1@S9.X]T3&=2R\UFNB/)L1]]D][NCVW2Y5.Q:
YH@3B6Z^U:L[b49OQVLf\dL\)-4+gBJH-Z.;2]L.#N?HX5PcUO7+N176=+Me0]:2
ES6BSTRLVS/Zd1;Cf]LV^0WM?fBX?H5ZVVV/4?JQ;8S2gc[d[^-c91(WUdZA&\3-
EfSAg#8ACdA@]3EKH@E\2>[P;V.QC&H7[fGOES>Q(/\GW3[FHYd@)Xg5:e74\GJB
(4>Q?KG]3HeLO#g4@G&BZ>GZ-^5Q6H5_S???f+FR,+22M8:2:d>W=8N3\>U;^YCC
<154+I-N8.e\7dHPI/MZ&7/5BB9XG1Pa]^^MI]VeCU+N6e.b<0V7MG6-5^LA9F9(
?7,+V_FI[g1LWOQO3/ENg6SX_]L>M]f,aZ4G&-</O0E.3ZC-B3\]HUXI.PaV#g58
;>_@a.g.4@Z_Uf5UYd-J[YA2TN3Vg+SCP=F_S?8HW;)c#IQMQ[da?CTR13I\+[a4
K[SQT8D7;=f-WffF@-1/B,W<eN.1VFVX&fe=6E(3?&1[LNHFc^W+OU.0<WZ_2]-Y
_WQcT5VGd@+#LbFW9<XMLCeb>L\-Rb1]e)O9\8;(85+1<82(5TRYUHJ5fC#eRgX1
L>;;Z;R;P-1\OSMCOG5(+3XQ,f3&J?a?:ecK@P,6RS@Y92-fBU-AP-4Y;1A35[g]
@K)PG-UW4NMe,&343/a@b=P==.+II7VT&7VI>L.@6)U4CFQC3A7dTM.c.C]2;U<M
^AJ(OJY4?#IE)fB5)LX(:g_N3+480D96>_F#H)FNecA^_77gf)#T#U2Z2c,G+6D=
3+JN<6D^4)/bJI?BDEL\7IQK_\O?324>DLX=Jf;E/=MY0F:VR;b[?UXRW>0-dc6\
-A2<XUe(g]NZ]4_]bagO:M53c>1^.YT@=C658/&C2.X@aUQfGdO&gVWYC])FMJdI
=-NVXEF#O75QNZ:G5-8bJ<E+OF1#ANa>F3L^EeR6eY6>VG7_@Rc(FEbdG>]:/XAK
N;f=9=YOP&7Y@=a7OKR74ecOeB-6NeWW-I;V1=(>>fEZ7>2.(O_V/;^8,<I,6dWK
&,6>b;U\[P0g8S)bD.T<_Fa-;GXGR?Z3,&1BJ_FV[c,]KWR>M;Y+0C3c=:b8/6W@
;7Ne4/bbd+E]8J[OP;f<d((XAH2g-Ja1IN[^QC>S,7eOJ@H_I^.V+3O+][e6AP2)
(Z9.?)@b/6N(OEH[g8VUec_U>VS9.-8>.0=F#<BP[=UWJ2869;1@H,3IOgJ;8cY]
::FD\SH9^=2L60Z_N0WA]\WC,,T?I,K84@L2#SHM9N(^2#K8CS?74QD:QCG#^(FB
U##ZDD.ZZ59E_#ELe=B5:d@BOMS]UL3NB_(S)]BZ1_,=LAMDf#[Z<TYY62e>Gg04
Pf>f[R(c]cKCB6Kg4+.c.(Y[/7[aPRYX-:5VWI?#Zbg/9V^/S5K_.Q4J_>.@NPG8
0]:,[[4M@)IS,2XG:&+U/c&fd61(.]L5<&:4-TLcV8Te&[B/fV;:/9Q)02#R1Ve9
Y4I/B7fSa)PKMJ#d:YegbGA=38A^gTF:3E>IIA1b2XK^PSQWFO&HA-8)<:GQ/PLT
OMQBJagO.M7aLA<H_ce&Nbe<OC&\UF8#eEW>\:I-&Fedf(1DCAK1<;>&g6CSQVWO
C[e;:b@FNY&UFG<P<BB1[g2OgZC.Y4,=AGBX#Ie7S#(QFX9A1KHWP8EVS)Yd63&3
N(=&CFQIX6#G(eX6aMX\^6KQLYT02/(Q2&ZOGGca@18ZKU#f1]Nf8L=9<a&EP4;?
d=8OLM8S:cXIF[[8/TWD5HFMHO:Y#@M@U&T@bdNKKZ[gf\(8PIR\E<21=dJ\LZ54
fMfa6LMU\M;7\&0B.a(c,+Ga]@>7PY9<f50dJ\ED4QYX5,,H@f[)/JGM/O6bP.QK
OFP2=P:63X#eUcW3((\(D.\=d;3dF+2X@=Q=Y/:bW[KAOE&PV/[ad\IP0b42e:QQ
UJCT-^,Xf#X0.DC,8?\/5,BF.25#N4[6aJ&\(CcPJP(FA#=N=ERHgM.XELUD:(;L
T4L&1b)3_^NH[bDG_(.8HSC7.g/=N>G19F]c9=G;(P0RZ>ZV&c6MRM;Y\;ISH_#E
CFOLZ\UG+TaNS[KKAYdUXJ^/V@<#NQJ6KX;]QQLD.@\+X.Z^d:EKMVeIR]Xb1JC2
_JJ6EB,C?UO.BNaXXNb/fPORS8.L^DXS)>@b.//,dKSG[2BL(Q^DNFMT:(f&a&=F
9=2EW\QCRNS;?[JZD5cb[H(5A==N&_Ge6=e^H[f;;AW&:&EOXY06f3Y_8N#ZZUP[
d0]+G@D[G(D=+>.1L32W=e;<_+HE(4EeATc-23\Y5bL\WXD]X-C+(@D(^:QS1,b<
C&-]##N68b;GF;gU\a6AE,+F5Lfb44bU&b_U+3X2-#(d26)Y_LYK>U>[\T>g6.IK
bPdLd0aI<PKZ;7_8b=eY2^>X<D^O)>Y3:bV(D(9G.[WV4IXc5KaM6Re\N;a/9c3(
KDAfM;d=bIAP@.Z?10#0M?NFgWOD1CD,25#<Af91OB=3R2QA.\fNe6W/Z@O/X?bH
&0B,8I3e1>_DB<#,G[+g4,\.QNg/:+NH\7O(W6MgTJA?b.RM1a,_XU13c&bWK/SN
bVN2(PZPbc@J#01FBIL,2-JaAc?GfO7Ne,dV=IZVHI[YO:VQ098P9Kc(]<P>-/Z1
:=5eRBe0BAQ<d,R9E5J.CD=(:D,Y)G^-^;F;>YZKB@X+Q5W89<[VI1N#57UZgBDR
.>66II:H[],X=18_9Z64+]CU58X]XJI^5HV^cTW85GW66OES\=J.+UcE&Ea9gK59
[_7T6\=DK?a))ff[=\eT_()=4NQBfIR6_^@+6aK@/9cdDP]\^]CaDP6-BC_&U6=2
F#;O=D=RE]Qd//)-P7.QC1ILdM-/VGH_c=0Bd0:9UAb((GFgBG7bE,T61+(:@GJK
_V?Z8&0bD2<T?]/:@A@W[G:)SAf]XG8Nb:-b.>bHA=H>FNfS&U,,[^=-E(ZD:2dL
Z+TE:Y9^=&Pe^dZQ#.T4JDL2EZTO<D.X,g0C>.V=<L;Ee.]N@(]ZUY>55UN2M:b;
OC4P)HN(TUYX0CBG()R#.dIV:<9T2X5U&T.dP.>FB8U/(?H&S6I.?D#5X1B&]d&/
N;Z(T7N^HG)>Y7T=/5)BdQ(KZZ)+WPD;T^CZ+96(X6@?aW9[><[1^JX3Q2fSUSbG
&AE,C)FbQEPJDC8&Z4Y?<:X9f?AA-bU=)--C^Z2e2<R30P-Y[RA#&SfF-5d2Z\fT
#W(6gf>?E3)3O.A>Ka@GUf,BL=QcB,,ge<Jf3LN\>bSdc\B_L<MG0Z)[gP;T,IV_
VU^+(cUKU88#F00<.&.aX<S9fW/8/]6g5-#RC-=Tb/7Bb2^ge+12O:c>QB(IQ]?^
A=fF1<>R[@,,c&\G&a^ZV2HU9/YM2Wea-IVLBKa<)bC<FH10DZc9?/2ID2MQC]&Z
CZa)#M<KA\cWA1?,Ff\fWfI3Y=EVT&c76AL5+6@>QQL6N608(5+8JY?3S-=U3\<S
EW&F=?\L6dY9JQa>+<2=)e&Qe#a_UBC@JUVY>/:BJ^WIE5MVUH2e4LN6A&NBRI];
bOSR46F[>:R;d^SXA5Jd\,A?7FO548I6GGT.0606SF6_;:/=KQ<3KMFK7KL8^A,a
LQW.W0b>5ADH]a^)O2FHd7)VdBCPA[6<0T&C)J?[V30S@(c?JaZ:8[^8)&4B>@:T
ZI[eX576-g\W\aJ6/[K)G11;15W8M(IV_71LN3V4ZP[aPO5:f4V76IOA9WV7DEfU
5XO3D-@<c8@P8M(L@>J(MI1E+D;&4gNOcO#bY2H)d,[7+1]JYC6;&MBgE&Z><M9P
X;X/A:S&P4HXfQ3P8]7#=.Z1JQFCCc68V+/aWNJGb<c>ad21f\]O.Te3=aK5P@HJ
>C6>#_Df-MYM?@ZO#?W.Nb)P\c0BX1<TGHU54EO2JEdPCWP5/g9#=Y6cDX4=^,_M
,BES0WNKEU:D41P:,Z[>/7]:W>=f,M@\/-<;J+DgT^#H:gVU]d,=OVL-a5?7RDaU
d2]5aFL_S#H+H)RdQO?=64;,E?I2;I8F@;<[Pa/:X:;(-#>5GYXPFBABb4P@cV0I
cX^5+)^5#Q5.03Fa3V0L?-K(9=4XN(Q7/Y5e:BMgb?N_&SM]7@DS-C16+Q;C#X<X
]/f]/:3E\\cX:RXUIg,/U9?eL+DHOUEUH,Q+&g^\:A3;T:TObYS._+:@M=N)@g\R
.&U/9dU+eH\A_@WC\bN]9AbXNQb6A6NOa1?N@.1/B?b=UgQJGVXa6XD:=C<YgbWI
7fI:+b4IfB6@9aPRDUI5a.Z_d/T4CKV3I62XaLbTX7Rc\HE)g-G<Ee#C]0QFKg<+
D?D:dA>b9I:eaMHY&,A6B(Z-5T-I4c_7dL>+1f#?)WR+,GQVa)SRB]L/9c<Z[Q._
+K/@>K-FQHI1SQfZ_Cd<P+)eJabHbd;Q[G=B5Wb_&W:^W>QL52\J]XSadJ8TJ^I=
TPOM[&HK]FYTa&NZL/.2T=(dF82b4aG<TG68Q2d)KQVN/L#H0De56P7+-1Meb5c,
\Wg3CJ;TaT\CN?&?1B&&MS3)[fWcN4eJ=,-;64Gc8D^]AL32SKA&5)K1#8-LF1BD
-1;a-bS^@4N[&]g5GE2VO1;/eX(JX+AX5K<bN(?INgJ4d]FOV;,BHS_WUaYX2K_H
C:RPNMG7/.dC9CWdfS;S3V_Xg#geLF0WH<U,WGYD1]O0CY_X<A\ZM2NdI7Z5dJRS
31P_]d37OA1;Q@3WCQF/=>[,c1c6;TK=V]-d<(=4V8_/?ec+5=;RdU/[cWf17ZAF
-AYDW,&,R--Pc>Fg[&=50c>5<A^c50OI/UX[SZJZ[JCJ\UK&NQ6ZH[I=fOWDE)Fc
6T1OHU0SIaM9<VBDI6#f]Y@]7/=JW@a,R:bW@[?[07\D/_d8Qc50gfW-?6\dF/HQ
K-1&R9^7LB5964f^=N(b_<8f(Z\V[E+;BX=I)MIN\MUIFY&&2N)AaT]-@=B9DU3,
S>gAQbVeaVE1Egc_)HC1dFV[^&9eJ2Wd[70Mb8@Q_(1G-N:CS+9<RZ.6D8<Te\I2
FOQVL=4G<>O^eBEM8\N[dUe)V9IeId/X8,Q([OC.;X\K>E290R9&TbF(11[dZV2T
_6W4;.R<5HQ6F4659<@YbL?\\[WZ)4gGW;N47?X-HdZAD.&6I2bN<8J?0eKfW\SS
.:-L6LF=S@f?^[?=Hcd33fSDO17MEKfW7>DUSbKKFE\RMf927QEP&O,[JEL-IT&C
[10I77C?^L3e=-GWN[;e(H&d.U_J;J&[Z^VL[;&b=)3WLA(9E^IY<MW,LBAR+]@G
04MP^aMB<b&DSRW6BK[9GfF4aJ_Y[MeZZ1dG,C-I^6[U.IPJ&fOQR9SaM1UdR=,3
D@^MYJ_F?#6)8)_P8RIJ>O=L\Bb._FCaA-(/bDEU[YCWf/8EA,9TgB\_;ZX(fR.g
H(If^LCA&TP9;Q)ZM-W/\4-73FO+18PU]5IgYebTf0<58-+_9T2_,&&I(UF]F7DH
]e\U^3Tg#0RKZe4?AXX5D2TQGH?WCMK,2,QVLcB9.:&MbK)Dg5LW4S]DQ,,V3Q5J
Z1-C=^I==C^IQCP/]G=S6YW_SCT@(aI(O<Q)Feb?6bMB8WIeZQ<[fc=]WgJO7/\Y
HN85c_gdg[N_Q(ROLB^WM2>]81I0X8S6;04\W,6Yfb#G]+QIc&(;UJP^8S4VC7;+
GR.L2F:2ZZS1ONO]C-b_4NM.TE[CG;Jg(9c4_Xc@QF8E0Qa@7#d;cOdFdMbAHM+6
,YX=c1&R&20KA^(MQ<Df.>:NYA;E>+KNAX_ND;3B.c+X4N;c:X4?Jg/.Y.5QLBZB
RVR=c1G_]Z;,#VW>FX&Y<L7.QUHJJ>?aFg9df[91bOH9Z#(TRc#CQ+RIX?PU^]J)
RTe@;(SUL#P)JX8:_W7X]:G/&O<S#OKX&E3]+&H,&\:8E?:/gI@Y1_;[.)>DWBM2
6c:@.[7)MY20UC#B?OWKI(@d7U1/_;]\M5eS1/^KVd>Y<Z<b&-A/c4C&(I36fSZC
EfMd3Z&[PNB\>I^YcG^?>6>+ENBQ&-fa8]Y()e8G8-5[K:WUKZ^56BX.R,NbYFOb
-^aKLV]+AF-IAV+8,JTGLXXUI^e1VGScFQ74.5F.#\T;d:ER8:#c5PJ-+b<bCaGg
bW_E)N5g^DT\fgO>7Q[\EW9.g@A0J?CJN7KeAXS4^>(+B/N=VWcDH5WDA7db=WM;
96HD++d6F;<#cESbIFSK290Z6=20P[1^Z]/X_[a+_X1@I+:U5;\D0GE#CC1,Jc,=
CZ)3GgDd;4X]>C2[)YH0;f<1SfbF?EKC,g1bDL(#+9-S<OQM6[eD/gAb7(+O>SQJ
+\SXH&)]I;IF4)NOW:?gT48[97?R.ZW[18DD/U^KfZ=Jc#O[&=34]&AI75LTWTK\
.U&]JSZ_V>[+Bb>2\P)EUe7K,,_=2@53>IKM\A/)\Q:,)cOO++[T).?>Z??#<_76
(aF@MeTcJYKJ118-/#gJd&H2Ra/ZB(-P5LFV:L#H;-((KXE-CK>YYDaaca7c_62S
9-a0\&bV]Z(G=)(VNfS:<b.]AWL7OCX0D4dR6d&26.RA1&2OFKTN4+Z;\fQF?OVV
<:^@I-/U-/3N2Ub?MY>OG2.Z^@+eLR>]EbQ3@]\@O;)&CTZY@(PU3LZGW^8=\O2K
SIB8V6WALOR0<b4;2M5^U#KC1YKDS?Q1bR#0Kb@@SA0GeS#@OaQUD@f_(.Nb?ULO
E8bXeLN0f\@ACKeV^9(2.;N04R?_YIf+LGQ8:4?R?e\CM7P+A4<F(8BML=44Q-Q?
6_^M9^CMJ^X/GBdFbVR>0WSL1C7L4<2-_&M#FF3>\^&:#AW)#<]f3++F4^T?N#KJ
(HGd=S;>4+EJO4U6-07>PRV55:A_P=&>MHEGa+^fO)D@M,@7aZ,HW5WF>7TaD;R6
.bU2?C3>4S>68;KG;NUUX(7fLd7B6#/N3EMK<J7TFM]?SSJfE(/_dL<JZ:SDBEA)
4G7(9P;L(&QK<Qef0e?ce4_?1],DJ0+H-E>I/a]+8XM[d?b<6LTS6H1,H>KHaD+_
^8\,f?+g7=FEEPAP.fS-=CW]M7f7Ad[2_bG5(;:E(C8#-I_TMdN:=R6PS-_\(Wc-
N6T7W^?<]XBRg-<Hd1^5,Q\aT+MTMO:cgX<C3\+e2XAG<bKeRLZdf>g6bbd^Q\3W
B&QYA=N-<DX9_U2:SWVX\/6#^,::4RECL@CD7>;UU-)MP.F8:T>NMN+Zb3+4(IW8
^S&_c@+HCZQG?R(9>O\T^3GW]/C]/e>@P&_#=^XYVLF73;7E++:^eC/>+YGQDIMF
+F7I5R@+J5Pg/CP/>.cB\AH<Kc.D4N.gd@dQCe+\^G+]^([]LZ+ce,CEP(I+UPE<
UU<&1QUS2@B.WS:+Cg;LLFCc=.dTbMT8FCXSYM[:7^@a.EMTAeDHJ<QG\?4TZPRU
+RB-fAYQLVg4965>Vf.[f->:=D0MI/YXXQa0V[6:<RPX)gX-4N_TL0W-dMc2U:K@
9IU:CGRL81-].8e+06gLH\:W]^N>I0XHaF3Vb5(V-STU]1d6<[(RMa#T8=<S9b?U
R;IO&c-WXE_P=FSJCIAf+F(,E0&Xb04/P];9J_G#a1/8VW=c[^OeWCFH-\H7A5#/
1OZf+AR9W@AFSc6./DE4d>(FFFMJG?2Y&+P^?dC;5d+K^f8(^-4QH7FI__BN@#NR
;ES>C>6ZDBAdE#:LfZ,R6aGbFQP5fPHN-M/If2L^,0(?P#P,#9G53N0HPYHBA,dA
IY>6KKZ?;e3(+Z]=M(\H3ceZN=8?VI3&9eg_.U7EEEWc)N)=AQRQHD[+.GX@ScBU
d0/5QTfD@[WH]NW5=2d3.<d[[=)5N\GJ58[QDJg6.)/[#XK)7fPQOK-NQAg_aBf<
E]J0])d]P>3_-3c0FZYKYVa\9?30>AJOY>QP3XgD?[:XNE5D@HT^;:40UW8YQ(EC
5MC8[bA_/;^[N]P:YP<C,Da+YbK&1APbXdTg.g+3XX]0Pga[MRFP:-Kg?],KZb67
):)X_7#-R8OO8U]O/\d#/Z07ga36fT5bYfBJ^cA\Z^\;&XX=9QKIXFd.R:ZT,7ZH
g>dCND94MVg78=b7,+<gOQ;O-VX3BV?K6/1I9:&E@1N5+>(4D?=/IJ,ATC]82gA(
P<0F.+1U03WE&2:KeIH/5A^:IWfAR7?RcabX4EcE-UH=6>)0IccPGFL=JeGD;\<<
GT,7L@Q<M>#FJSc#)(NG2^)08JMFNM)NHN5^>U4bX.4Ec.:&Z)Oa,^Nc9GH>((F=
NACaaW1H98YZHP\;#47633L94D4>#dTAR2\O;&D#K,WTQJSYEfN&>0Te&:ac)V7c
Y,N2UL8#b.D_YDafG+ZLcVT3)\N]d;g(CK-LEbKfA^Y.IF<;APWT5b\D4e@@54HP
X:B+T<a#0AX&f8C_MAVW_Vd(1=YL6R]<0#T:4[I@O:^+FPP>^DRX+L0<#&CX8W[(
+2>2WVNfIdgNU&]O]0EeaeeEBd@BQZe3P]8c@/J_[IU)4_6#H,W,.^.f&(SIDV\I
/c]O8bc7)Q;VEV@H5a&7<L6\:C-A513M?#G:a\c4EF6&9/DbHNSC,=gK7A8B2PD/
;eA-Y/-ESE^K&H.VS3J2Z3IIcV+6+<\@b.HR+,W@@[D7UW]D-C:KGcf]=_QAc@GD
_DG-7#QJ_U9-,7Gd4[22SbK31bagW+:)5I3]\U81IH\VgIe5;3+\FfMK+NEQJL#?
/(@a4RB6ZZ_g6[4&YXC;P_@;33UFZA0a>Q-,fX5Wa1/5QF?Ma&N;-a5_DG@B2bU@
.(STW9\?KA,/M_)JT[BJgRBM_&,CdY<9./IG<a3HDG9H/-@FHEV=9?3+;^@F14LQ
(S:P/]b@DaUTP3K.0AfbUT&/UdEP#86:6A?)EO^V/fO?SYg@[L,c5NcAgL--1\B6
)P<U#\T)+62CF+6A^DC&LGH<GKb5-QC7KR:]2@><6LaAZ6\gc8\Qb/1&R/)XeMBd
>XYZR@+<We+0b@g-83;d]R/L,-15L4LC28NF_QF>S2@P&cI2W@Rd;d0GAb.,+M;0
-\QE]R9;L)2J8fM19-T@e3[IR#BJD>7]?GO/cNA<)NBQ[Jc);MM^^VUZZ#R20N+H
9FGDc;4Q>^eJ]gc@fOa@U>>(-5.PGbL_cZ:TSYS]_\TfN]96Hg?eC/M_^V.8+cXa
(ELEDVCaI[UIY4S(^60<T\GMJQFAM+\OfP8IWb#6_@8=)A.2#ELQ0.M2C.c7BSKe
YKQEO>^7,YaNJQ.[N6YefHD?f>I7fPG,g<U=:O8>3:<BY^Vd\?8a]7/b1gL2O43;
)gN6YWKTFdGQF71XN9/)f(H?UM-Qb>eNa[L/g<:V/@,+U&8WN^V75EDSX4XRB9g]
S5U3DF<,gTYOUN\YJ^B-e]c=ZU.X)6Q.)2f&P+:T/PNKN9??<@LRA(7^K?FD;O#I
40FUK&TR&S(R6FU<#T:9?KQaBYSFB6B3-=:C71)#0?cFg/SI);O]CRZbD_ZTSG]f
,&=TAH);E,[ZORGEfc8NE(E>\J\/X.6ZV=:GQ/V/3aH2J&<=A4L9cNV7,[f=.6=1
T(+/U1<U7a0>?:OL;:P^V#M,X.=/4HeR6[1K.QL6X<T+A@;XRO)M,3Z[dT:,Lf>M
FY\4Hb/032E^e)(d:V6&GNC.V];gY<@)V@F@W(,U#c2?AIJ/IXeJ)C64JZbLAE4.
a8f=YRea+3KZb>#(GSf^1TBLa7-(+\.1DT<F+KYbJW5]g]Y0Dc(M-T3c/(7)#5B6
9&?/T[4/M-d1g0O[]N@Vc<FX49M\M5\,8f8^^-d3CN+]OX7G+5W=TZd-?8c>\QU>
DcW3P.?[KAM1@gD)SUaf:LB8Wc21WM)e.Xb]YW2#AXUYC(8.^1a0]21G,Ufe29M6
EBZTb6g49e<_9KAO::@X^Og76(3a=:a2SX-GTC]&(>T&H>7dE_YB[ZP/C?gMMB[^
>0?6C/-6)@CYOOVe7^Vb(];4SK^&(M+I=408YGcZ1RR=D(A9;^9ENUPDL&RYA_9K
4S;A>E,#Q6;HYgS3+Bd?,Mc-[<]XbC#U_@BPD;AL2X0;45)dILfJ51JJeC19CcdA
:6YC5K8X<_/39AE:5b5N_CdEX+JE6,RW^&>.A@.4(:W0;;\3&K\RU\,S.ZCAc511
>U\]8&:eUN&c<?JQ)9\#L/YGU8D^_4X+:f3+/_8Qa6/;=,__JSVG&EB#F.D-g@8H
5a[+(CQ9D0;P\FW]\A7dKQdV,DJ+(2;4aH7]d=E^A4(:CFU81OXg?5Z:g3)@7_fI
3++3QP7YVT&==-&-f^QEb+>A?WE]dcY^[I9Dg3\I/I;/(\.BBO?802/OH,e<QF06
_HH+cR<D)fV99QI+?GL[&bN>(O[H(#6CKcQS4;KI1;>bZ=2^<Z1ED\3T[V-0FU+a
U8ST9.IG(4FKX2-O8]HLLDP2RB(A2b13(=(,IN\EZ&(VFN/I\<9S<GNFT&]dXd[_
0Mb:TQU)GX+]:)HDVc0eR-+T-cZTFe.CbURR_E>9:W<ag>_9R:#QLPdEa813./&@
f?DT2aMC3TYWB<L&URgR,]1OA2RQ;6,<9g/?/Z&[,:T&&UU=5MU61OfQ&P<eQJ4M
@(3>7JgR9,VFNH/g.NIU7\3/N)_2MW#gT(QEV6[<6K0KOF:(P4VB=aI9O@(^gM/(
ddgPGeC4^E(;ZeQ(76cOU-J\/e4?=KT;Y;GAN6dF3K5Ke5]J=[d#Z^7S=c@QY2gY
O[.T?^&7DQD#XZ^ZM:W;V,\0.1F/V/KHFe.d4f6#@WgWd[S6&]_BT\9bgH,8Ua;)
0#.-c^W8bHFG=OEg[NYL_(Z6gGg_>0:(HdD,KK@2WcNeI^(K<::De=1=Y#IBBda8
]3_X\4[W2GddNf71:@EJ-0H^XIDNFff)X-eGN83C3;(_^\)Vb-V<OUQ;Oa]A7@5C
18;eE[=FTT@IRNN_#//f,4@@LY)6J=U8L-L&+0TB&F-b\>I7_.QE^\^=[Pf;?WHd
BdP-A^Xf]e+gBe]f6HOHY;[S2PFQ,/g.a78d/KZ8WZE-B5D#dcI9#GIPHO3@136+
.TbT/#NEa;]X(/gP/3\PHZG13f)=E?YT&9=HeYGUe]H=M&EB+X#(PVeSOda]b;\=
<U7LQLeg(@;A9aM[J&dU/2CBOA2T9XCO7W@Z6F/R5>=Sg1L4D5Qa295SCd&0P<Lc
@X:/=-&EQV#&3I(F?Y7,7+5753LSSFFVEZgg2=MGa@XC=29E?:]\IEU6/R:[KWAS
cTaR,ZaCY7(/D^U-g)A7S.TVTTH/Z\8a6a];<3=dVGO0Gcd@_d?c#+X2Oa(dM^1Q
V\UT4RaGD=C36M<KS>,dB.Zf0SDEZEVN>?11DQ&OB5f+94:S@4JHO1@AL#?PL:WN
8QXgE9dU5/)\MN?9KEZA_R;;\IC:B5@Y;dd(X.W?W]XT]EggM2)_LSG_U3ab:(JI
XXX;MF@KdN3LO^[LE8J3D,0GC:S2DgO^CFTSVfgZIS.@1>C0]NP#^M#)T(PDc\/U
e6/^AV.&1/5Q-MS0?aL&4WK)<7-T9f</A1M9\BIbNBV[a-0_c\^P4]G7_TR6)H3F
E]b2SfB#UU=PHP#]89(VP,+JX<5TMT+B)J\Q@Da25HA(e/d:\[@/@1Tf/4EC>2@A
/#A8L,>?FU8:SQH2W54]c^Y&P\A^d^cVT@6YW;_b.[/4YfQ(8O,Kc)Y4_U2Ped@:
85FO\-JAc/\B+2WbOfP3SWaOWP^@W>45(?2b:a8L<PEO2e),(SZ3TU,-).4f,]7W
BI(UMSD/fC)VDdI0B3a_PX<F@OOMPDX7(\)gSH^3Nd1<M1]EDR:\2XB1<b4]#.0M
TTXEMJ&^-6+;R>=/6V7B<O(ACTK/4=>,[@Gg+Lg-IIW7Z+)[W=Y2]#T]HVG]e#b\
JGWg+EY8>HHQ9]KEL#MFO_^aQU/K@CW>O#KJS4K>F>DX.6Tb4B+(]3LEW_gdR:0+
]b\K/d8NED+\eD3d3OY.X6KL3ee(2IZf.P]&#9VU;@QYUb>>#)5<#W8::A-(f0BS
7P6^.aEGV#Hc#P#VELK[:\74#dR=/S9DLf_=(GWTU7VA=36,Q<dSU[6)O\\IKTAI
TZ.PM=&,UZP7F&aQ4S=cSe^Y@X_Y^1Df_+OC6F/d\<A-E6cI95D9QB[XH>]S#2U?
Sb[gOg\SB_MDR+HfD7=IE<DSP4A?]+]a#/UV#A\)=\[UG3MIMY1<J+c;9N7e;OI#
3G5f#T0N@JRa=6dJ9:WY]3<?>YRW>>g2)#V7+:Z&I^CTeU6&CL/+Q)H#;2Q5.gBZ
+FNGBScA)-efAXOeI]bNIf86bCR06F#[<NFf:&dFd]G(M(Z](CG56[[dQH?:L?Y1
^e3fQJP60Wbf=KR/DA=KMbUEg3e7MLS[WWZdS[+Wg,3_[Q0-J.0#:6U<XI<RcEf#
V72XFCHRU8]\6FHc;W2b,Z=V/+Yc6F?e..Z1S1WJ-cR.,4]YgO5D4PMUM\-+20E5
_W#]<fYNMJNX0c5:Pc?#TV-2_Ca-d>Ca6X/?&.I^<9fbS6)[(A/dHH?NM>c#VUcY
[&^DagI]7f?EK.53,+,5eT:3.LbLeT?;7<)@3[\JN:,JV:A>KP@2(-:==P/a&;_6
>bI_g=d@781D6R;21,6-B(&)(X#2375@V?Me^AXR^4)Q:KPB_Re3RV3/@@>G&beQ
36XX<270b;7.CA,<_)=DCV\_+4<D\]O]29.=L;N4FT1dQ6=_@]0G?F&@Z3RL36::
Hc51NIBeF?-1[&GLS3gD=/D.=-,c=M4feC<L02)5+02:B[-fb2b(^THU5g&7?P^)
#-?;GBT5H]I=MO+&((-DRdOCM]W=N[9Z.YD6d1\#AETQ?<R,EE_c[<^P0R,9YeG1
H3b_J/0@6T1D@dJ3P#Lfe?:)7)K<fM:HPAE[Oe=UM_3::C(J-DW61L0dgVTRC;7d
=79/GF_a_V];^HLC,P_.Udb_74FAF3#TKR+-?\OGA<5J;H76^BKc@/M((^:DD(FA
OWe07)/L^bCLH;#(1N3VXNaMU>NX9aO[A(4:R2).[TY<C]6e]>]b[UQY),TIQg>C
LS=ZHBSCdAB/>Ndd/N#Z-be(Va5KcY:H4A0&J_;M_c(:V];G(HMeDFbRC([<>-(5
ef1Fga4.7aX_J[JLgCPSDM@RR]bH3&OaNb_8Pg?[6XEYgg8,;gR.J@TSPX9?,XPJ
,;)^Dg:X-]QC02&J?]F;-;\9_3<B,?d<8D6Zbb2B)J&>OX1^@64=A7J?ZIg_c,De
IH#a]UJ#WGJK8:8d[Da?62HLEcD<f?8NQX38(IgM&PX,,<g\]0WS(QFR0_ffUYE-
#4\>^W//&d+J6\)N:H/V2HV_AB]WJbJ)(>0:QbbZX\84Ob-956eP-8PfgS;SI46+
-FK<NH),T)b<LUdfa0;Q4cL#A^JR^=-IG.T80SJdJXVR8NS4[#6?7Yg#-DSf8^W4
X-.)M+d-4,_OK=b(;;15/1b<9fYG47ZH,E]W2WYb;8H6-[S@6e&-0=c5M06Yd>Bd
Af:,C.U3LXFR4?GPO3:7G2E46N&)@DM5_HN9Nc7d2HT^\aST:Q]4ba2T=75Q9AN3
=B/3G_FB<_(A6cQ7JX40;b:4dXfI91?;9G0V833FS(I/WeMI_>TfUbQfSN,3_0ZK
(VK:T?I?G^/9M7&#<O0)FH2-TV_/#K4Hc8]D^10Y+B)28=61NJA2S\YLc^LR:JAG
f8EGO-UDgZ18b:g[Ie#(]d-JG1@AgM/GDf+@gB8.J-#.L++DPYa1;B)(3)7/.Sb)
3V2[/B>V7g#e.?d8>&821Rbe3B6d7_aH14[#1E-g(Y+DeTg&Y&@-RH;)a4B=G/Pb
?@BFY;X=HEdIHBV/gEe,H8)@X,2_<&H+GJN&c<AJ(?8d&U:#(4:-MWP-YIK\.PO4
(;fZL/?#-3-WYOg<Q6fY>=L.1Y;<;D##7,LKdcE;bVeJ5C-Q98>(WCEg#(H2)-\f
92(7bc_U0ARgD1CdRA)>A.bUg9AfZUY_>/6E1NdV)3NODH7@\/<9Kc#a>:6cf0ZQ
L,&_Pf5Rf^N8?WJaR=EMf@#9#Q@@Ag\A30\eI9b^PN>][</R@T5_2<AZF3NURR+Q
T\D8e_:JJSR^5/H?7LQZIJ#673Ud[STB]6d5=H5fdX^?b,,;fK32>\3O=A\<,8D9
?[\KLXWJ<G#PZAE7K]g#]-G4f]@]<9XH:cQ:1F:K[9?GN5e(RNJefI--Va<6PZZ)
)N8M?>(T2CVU&g]\]1LgP.IR-G5>FW;Y[Z4BVQQ66B;:.UT,F?9G,aTU:Da;\_C5
[#?PLB1(V,f>aGWXV+7aS,?6](I,TQT:b]78IICDHYT5,3MfF>UG<YFJ8BEK2RS_
FWH7<B>KDB8AR[2AXAb&_9:+<ML/BY@DYdCALCD)2>FIPT,0V?.A1f:E95b+?]+W
aX/?+V@HgUd7\-Y7>WO9X2.d460FTV\E)R5-6+9^(V[,G1CX8=X\X^^8)1</Q(:Z
[7daB6B/BB6aI[,aN>,YSQ1@TDH@61Q>E3#FbI6=&fI]U1Pa3FSR5F96[)/)M^JQ
^B7C@84@ZA#(E?,@8T@5>MYJ&[fUf?RR[DJXb?ZKZJJ.]QDJXD,&G.7XEQBUTCdS
SNIQ4dID>IVdYKcPH,W/W+?;,X:CcOYP;^AL1^Zb?]SP&JJTG6?Hf3-6C@O^]YIY
DGG_B[/Ea[CT/D)P@WTY=05HRgeJX;#Oc_:geQf(d4N;P&+4f(CT425XT_JY/2MV
.)HT(<I-JSMXDg:VMNE[YgRJ7JHGU6geAc[PJc.cV&HgD9,d455XYB,c]:;?Rd#M
RW+GH@cLf/,dc+#WTL)@^C2+]2CB,gRNHVDTC@g.a^fg#XF3Qe@9/K=1\T2E9R?X
9c0^Va-IL7)DU8H<ddbZ]7<W9fe@b.bGaH#J)@UT<Ka/0d2PYG=4d<.6,VCF(bJ9
B]:KGgaUFT.CV/833XOcaN8;7PWU5b\](d[c8GJQ0N[D:8&UTd5Dd&K38=_R9b&0
(^KbaTB1&GYcH8.dBGX=XS?E@0Md=]@8>Y>Z>R7-V>)Y)\NAcJFc8c-Afe7]Y()e
d4XTP10VFdSJM@GC85S3]XB9-Z#W[a3Q_,G4=3C5:B,(gB+/G_<5ZPG;/gRTQ3XL
4405D0.cM_LeT[ZD\)].P,,_TGa_LT;\A\K&6OS2EX);dW;>fG,;/).G(\&&4-d4
;O)1&W\0d_TO^NI^)L@bXD6Q=3++2986U>-I#DG>g/YEM2?Qa4B@EbW:77+9bTLZ
c7BS;0ASJ/<8g?R9SPZ>0/PgL3GVLb>,N<aKD&FM147f^DcAQ+S@G)KY;LTGYW:M
P8&R1_4cDA<Vg^,W0+a5(-UXISO;P#6U,\M.J9Q:C[+S&4Rf1ge>;IFa(;.ZX5Y)
&VaK\;.TfSC<ZT,8-2I-E:,S)4Y3>b75V,R,G.\219<dTOZ2g,RFENYcf(gXf9#(
BEWe?YIMC5=YVfC:YNA2+c[/_SgZOJV(+fD&I7XI.eUZ(]Ka.G.7BLQc<VGCM+PE
JUMOHF&K+I_O:8GO,8Z.YWO?-+[X4OS2(ccfTEcZWBL\Zd:9,+(?2=AK[9b97XaQ
WS:d>@2f<T7/P\C7X+,B85#(L3Q;.LU(-e&JP;/\5<6Q+bMg37:WUTV#UH#=/=+/
Z0cI>0J07T]-VS>A?IY+\0]Tg+HGQ;\BIKEGOeRP>d(BM8,G,Bg@=#UG=AVQgB:9
(BU]VafG;__K-MA;1]?/CHWd0M5gOg5Q)&AX#B:/IUf9^TW&O[)2PC6[.MA;,fO:
Z:YIEE\OGHKF9:fa.I,g#1V_-B.RRI/5&<RIN7WO)2_S0OBVTbFWOO-_^c41O,8X
cF&]3gGN?;+<+H5,:CHAK+\H9,aS)E1-=_Q.W0Q3FIWAd?4.E_bCJBM\]G]1#6(\
GZUgQQc:=_BSW8ZQRNM4=SD@Q\1[P]/KeGf\6]HUP4Y1SI[-ML@Y):BWUO<?ZS1g
MdG\cU2#NG:a1H5R,@G^6MdD-gZ@RV,FAGMS.X&HV3g3(V4;1G[J0-CRDDTIL=9f
5NZaLY96=@^Scae-<:V\M+]aB<&7L?2[,Z+:5@P7F<&9aSA,@fbRgY?+X,/=&OY-
QXT]FHOE:F.MA2J0,C4;c&)>Q:GdJ+-HL^P#f(=De-WK5A+1Hd#D6O@53.(R.VKZ
ZS2C[GY8;9?CdA<OP?DQ#S6QAI/bBJVdK=DB/fGHEHB_faC.d;>g3dA0c6[<+<G3
,.FR&gSd-g8X3b[LVDcW2N<#;^<?H;#V@I=TEag[^YPbFX9:]20QW6:SH(c4GJH#
]17G2T/(PA.]LU:@(0#>B.=)[^JK&0R4/[\(E)W9+_M2]fFVeg,).7,2U#)P5fQ8
_eG#>T&TOT;LN=1Z>F8O5S0Zg]S=3gV&,L2H+&N:V[[QK_f)@R3Zg/-1XDPFV6T]
E6H,_9ZeC_fcPdR8/T@dXTU]W8b)PCLA[1]-?Gge2RDZPP@8cIP+<BY9M#;#]OIe
5F8SNJ^;aI<\0PLFL;HOD5?QQ3-PX7Z>NM@]/O>]HY^FJ0=P-P9aG<<f3]N.,-QE
788:e[K=P@WYa9e[HI&9CFD\GZL>2cH@V].A,WARYF(\5SB+T4&.]I3gf>=V#?a3
0CIJXK7D^#;P0I_I8-W7@VU)J(W<@VOPFBQI6de)]^EecL5S?-X3WMC<GT32RIaH
2\0+87JE<Tgd6D&bcXI@QI>>L;bbQ</cS9=BfN+O)&O=Fa(?X8g@-e8J\PADLc8Z
Oa&NE;A(&6IJ[LY\a)7Y&4<)aPRSQ[Y8D=NRY=A,@ag.L[\c/Ybd7e,S:&-gL@.=
_U29MAALM_;OQJR[>5XYC6&Oa58#d>3H&DZ0g<fSV&Q7J?bM]MZ?O1)W:6WOUSZ:
_4HH8.HK7)7BfeUS@f.?ggZOMH:MSC;XPbPaKI1<66^U\#&5:0N+.:K<+8aHe[_;
a.#e,B&@60S25L4>QFBb1H]P;Xea\_C/PW_Tag1-P>ZRCA[NaXI3@65<[IW#5ELa
3V::/\dAb))M(IDWXMJN46b^;51FL3YM+BK(16XWY\:dP&EXdHV_Yg(IG5LN:2Qb
NR78RBLa+LAfc0<=<<cH]IX7,2U6(_QEf(#Z#;\Hf(f.KTJ;VX[JdR?JH_<FSK+O
Q,=F9bYU^\0dUJEX6V5MUIVND3SZ3f7TWGNTEcdLXFJ\d:LdM92A#DcEN7[<4P[S
DNT2LWcYe:5+5]>FA.:SO=)/Ga<&(TS3T6LF@:PLX&.&@dg0aJdC?RZ6OGGEgF2[
R-,\4D?bK?;\WUU1Y<TSK^3eaMD)J87>KVA64g/-MQ@;We5=0J>@BF3c,+EeU>D]
X8XWa\cU1G#3SP5@])-=fJJW.dJ_aII4^(dN4QY\A)V6[009-<#F#>O.RJ-Z1e#Y
eVgUJ,++A&?4e#GO[a@EEV==CJA]+Z20-&BIEd+=U@D/L-.I:Zc3IS?3gM&.1=\[
U[M7/aBb-]8Z9<SR8)G-;DC0QJRTGKbe-6M5QMa\ZL/>Wc+-c8)C3=_X]^8W,5<#
8Z0=L>-<-HN8[(?1>77#Ed)7[K_U_d\LA(Z8Pa.7e>S_;8>R10E#_09K?-86(-H7
B#P_ae\A7a,P]=R>Y\@Q5>)76$
`endprotected
endmodule
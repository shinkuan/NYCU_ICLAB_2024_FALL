
`ifdef DRAM_PAT1
    `define DRAM_PAT "../00_TESTBED/DRAM/dram1.dat"
`elsif DRAM_PAT2
    `define DRAM_PAT "../00_TESTBED/DRAM/dram2.dat"
`elsif DRAM_PAT3
    `define DRAM_PAT "../00_TESTBED/DRAM/dram0.dat"
`else
    `define DRAM_PAT "../00_TESTBED/DRAM/dram3.dat"
`endif

`ifdef RTL
    `define CYCLE_TIME 3.0
`elsif GATE
    `ifndef CYCLE_TIME
        `define CYCLE_TIME 3.0
    `endif
`else
    `define CYCLE_TIME 3.0
`endif

`include "../00_TESTBED/pseudo_DRAM.v"

module PATTERN(
    // Input Signals
    clk,
    rst_n,
    in_valid,
    in_pic_no,
    in_mode,
    in_ratio_mode,
    out_valid,
    out_data
);


`protected
Mb&OQC0f-F6V6DgU/VQ2W&9Ob-,#I.#6MKOg&ULL^)(_8/c\YJ:7+)Ve/JCN^SE_
(J1MCTW[;LdEHY>af\R4f&\?.4P[T>C+@$
`endprotected
output reg        clk, rst_n;
output reg        in_valid;

output reg [3:0] in_pic_no;
output reg [1:0] in_mode;
output reg [1:0] in_ratio_mode;

input out_valid;
input [7:0] out_data;


`protected
EC19b<\_9.TB_>^d:b#0KZg?O9-Q07a?75BY=Z-7(Q66KMW&O8\+7)5?VS.7/[a6
GD68ME5JUU/79OL@EUaZcEA/G]M_.Q>]96Wg^&M8HMI.5-)0HVRdGaM,9\8BYdb0
be[O+,FSafES):T<>]OJTHa=gW.#NK4FY^_<&)2]aM#=;0(R,(-gG)=e2g4\?c2&
eE^BQRB0g/eLZHfS2YAXLV(7F[bdOFYbOg+?FAV,66L\+V90FaeCQO?EdPSR0#>/
0L/;@+Eg7d<<EFBO<b@[Qd;\-N^DQfOFZ35W>;fKYW&H]1R7\fIO--BBY^5JU9X;
DcS0G6DT0[0MBPAAZ\]>JF7U:N9UaOXB2]I[gP_/)9N4YRQc6e\W/9^CJIKBRKXT
\V-/A;N7)U_B0(+CbRBN-<,\HC&-(EG@_1Y;HbBB@.()U=9QAN]V;+e3UEZgX&;D
aa-)Ce4FP[\:QD/TO_4,C,A@O#9X:fd@==DPCcBD=0#Uc13Me<W@/AN@.Z:1&@2d
a<SgFEd?e_)Yg<d:.#K-c[HM=AaT0:g=e5R_,eIHC_R\^_M[SB_LQ;^TfX0eCCGa
\0AX?<,6bHaJ;N<ITP(?J==GC#P8-ZZQ\eL<HGPg3c1+ZNBg07J@<&<>.)@INc>>
D>;A0gIBSdYC;59[Bd#]\A<YA/d[GGIPSZ>-TMRZ6U>HOV^6TQ7_6-7aSS_+QH-Y
@eNQI=2fZ:2E_[Y4X2dM.N<[FbB02WgF_-@g7:MLV.W[U\ag/<YM>.(JC#V=UY9d
b40YdJ<=\HHHN#[C63?5>@&-3g.eW?[;DW278A-NI3,?;/8W\<fb_RWeeM&GQX8E
W)+H6@(\T+FU/]eOZL5^Q35_HS<98T,;O>0d:X1OeBg/N?gbFG^6H??-7,2QJB<E
,<S0W>D)KNKR^/<@_g1\Wa/L^X@gG59K5=#e(?J[g@3P3e48G+7f;<)812PNLDW(
NEQ;);.UX-#\]UOI,V@=B)E(NO&3,IN6FHQRZO\AJD-NCP[G^O04:3HF0#;LcbgB
2/f[H9f\BZ/V+H3Y\d(5TIGPT,;?/B75.&0&bCQ/N_eYE;T(:STcVeQ=5>&[S^8@
c40;g;Y2I:gK^)PP2CFcJ_0DbU@K=dDGS^R/YRcTffGP?M:E]JYUMSTCO.MP0,7M
>3[e&D49Qe]8[8M^AML0KN.EHJT5d6<LXYJ5C-,U1TR,SAK0OD,aQa\(T14CVgGT
?JJ/_[]Bg,\VDa30<^c&<-gE\3I-32MNA.:,+QW-_a+OfWMUXZ9,<7:a@Z06QP>I
DNfg-IC]\S,f^Zb54XM&gXdWZOMET8f+[\D]1BJg+KU_&Pe4,6D5G];/Me(b1)8J
@[KE8]1G>=1S+H@b2FK;00dAP.3P;MKbeLURCYA?T+YY\f6T+7-faIf@D1HM8F8.
>RaLMH@)c:1LJcY;:e@g4(F1Od<0^/A7U+S@YHBdSa&\OYbF(@Cg&\#R28B7F^1P
G/S02b?eN6T^GH0B,c>)]LEe\LJK)9XXB,E=bO;Y&^=gc207Q\Uab3Vb1&BaV1K=
J:#:Y(M??5P8eWe1:KNC@IP]aUaLH:C])@K\\/(V[43,RcaPbXMIZ;W#5Dc7POMT
G\]G;D=?QOCIa4S@aC(gZO7+N5&IG#fUR<6Y1>Rc:V9PLB@Gd7gR\aD:.SBAZ)>6
:0#bGG,#8;AUdc5RY_P=R+X;EOXZCJ=f[]P6)=+]bCFJH8Z,?+fC0JH.?NfU2/Yf
(DLCZPOT^WI6fQ)AB\.E:TK,4;FJ16M&g/Pf/^FJc2FAf,6)g/-Z-@V5&aW8#44d
+,?U86G1/]NdL&HZ:(MD-2#0=:_gF.(6>YN7Q8^(1?1?CHKHE2gON[O&Q,\RS/<[
+\:\DDM-9DQ@WUB.MAfY\)JeEBDW1F=XFg9eBe#_]G8U\CU2<WReUC(^Bd=@F:R)
VB53PTeXe)GHU^<X(aT9I04EgZ,8SCZOWFV]:,<6)D_g#bb7+EZ;_;HST)WXUQA3
.LdccOC5EE2(T7TbTI]<SH>Lf#+<N@A,WNPY>D_g0K]f.Wa3;O&Zc:dVOD7OB)4Z
V24VSR^?H5P2C^)[f(DAOd)gR98/15S_:b@eU+WUB4B?32d3;(=]BW[B_d3AHH/J
ANMG;c4\4[0,3R6d_]BcPCBf)5,cG)43aRQ]4\?QK9BAZ\e<fP/:SIR);PN/F,_[
^NJXg):D@U+OZ9SQ<X.AXK92K:F3K3gEP=Ha.@/FD>RZ+aFX7?GDDgXR/PQZQS1]
XFD5bA&5[[KJT,>_#5RFV\]LS)J&GIb26d/H5gM:6c=GgC06DS7P^4\;?5a-IXSQ
H/:c:^<C>#FO9M=SaT<bU:G6314,K@cX(+AV13IXS0UN:E;ZEb?,dD2cG]_[3VfY
Sb\XHEA8d2[Q:/HD3(1)^d0G^]JUJB_]Wb2fg;Jc<VRT#=&beE,X4?Ug]=K#EYb<
VBN&MVX3Q36L.,4CfXW^(8=.Z,&3,.EEJ@.L@X/Vd<8(L)A&D<2GL.QKE9gO[;UQ
V\,/YUdF^S&+_cg+faC:3Ea3PS?5(:^.OQP3XP3U3.S_.)Q@D@7IcTGV3^Y9=eDT
,(BJ+W-7&3g6&[F(JL_X7Z7Y;=[KY^+>>U?2#RS#CR1PCY7C1IVEWBO5X/:_Y<:;
.=-V:\;N):^\Y3R,gS_6TPW:F,dW;6RB-W&_</IZe7);DefG],7<3f.dZ&_b]CU7
ZG3,@YQ9FO?::7EdA;fV3Xg-1eHfP[D#QQ6cHH9SR;EZ\Z+^2?V)6bQcbK@bb5W@
;8>KdPO,=XF<?::SI8g_N.Tg4)G.81<dE#56E=FD+>?++N8CK\5>_PP]98FA;/2=
-LFF3H8;MJTP7fI.4:<0_UG#Y-DN,O42FD>3J#8#9X=+EZ9Z,gQfgc3VK0JD,>WJ
2W>?+W<Y6&0K>GVRHO2SD1Y0^Q)_6V+4./1)1N2gJ3T6:;<2>>a;6Z4/P<(1_+F@
?a^1fX8&eKe@YPL3T@gTD<^(a9P;6>A=ZBafWa5Za[RZGU[WO/S[aE&7\fAX_f86
g_Vc=)^A-=VN13?]MfOC+J[[_8FX?XX2Z7OE/NgTV@g5_3JUc.;B<I+fGN[Ga45,
DeV3U^4XXWKB@=0G;40ee7D(+=B@>COW.Q4I1):ICSH4RMK+6A=TG/72.<bJLI,/
-8<[/W:gI?HYDW<EZ_9NBCH\J(g7D)L\-0&.^C5D_?Y-=CM(;U<0VG9?,]/:DZ3/
V/c&b?=gKg]S9WGO7&-Vd@(R>@V<.Ud01^?S#3[eQeB&Be>[..-__.^3#AdZ)HIF
Z=EQE^#c;cOLMFTGB7UG391YB,##_dE3<DUcdZ_6,d[VW;Q?SCCV(=CF2LTgYR8.
^DN(Y^GUd^?AZ1#aJMSPbD-610&G/T>(^P44P+U>X_K;beG9SYGHdfC=WW4Z=Y^9
B[]b5V+&:g#c14dGFE223^cYNN&-R3RFUX?@YE.]D;1c/[aT:6eAZ?W6FS,2Yd(M
N,85)CK?E2#gA0_dWaaPA]0#2)/3ESL(-U+-1>2,(b[IJ,X\@B&K#TbA4QXR_4cO
L-QcQ<+9#F\e6:R/X/(PdegOW]G<GO;1QYb1^7UKJcgU/OSLfbVD+f@c;/Bb]G.0
OJU-dD]b2GTZ\2RUD@O^TB&^MW&J20Vd4Bgc7+f8YY#X:0X9=b\L?)[OLVf:aMIc
@I1-E/F_fF[XKEMHd-DNcYG.Y[@E1/2KINe6;Y063,MM[W/9E7bB52B/ddd.(\:>
Ic9=<S2LT?5,#SR0d[?7YI9=C5O6L9?&M=fV_C.7T=QGW))N?HL/9@D?@@CZ0,0+
CI,Z5T9cDa9/A^1]LIF\<B\SD8]E0daeJPLKAN=\;3?SPBWH^<3@/g<7-dB7S(-O
GXRPMK,Vd93ON/U]?QB,PZG#b,6PRWe\?b.)[61H>7XR/-5+Q7G+#;f09YeEEN,e
/D9=YQ\5Vf]-3g[V.+5QPe6cCI&3cZ:O+5W.HN/b4AHK7U3PDO.aAH\Jd;CQOJH[
+Q.VM)HA9E\d[RC-SeS\\7WR1719<](#Z5;@XB&LP,0U[UY<>S1BLUJP4.f?L8-?
;)>QLe:NH5F\Y3g?0IE0/P,\OZ+]f)_XFbbU&HPIDYZK)69IE:1gV830LR5.Q-N(
,VN/e_2[ES2eE1\B.Y9GFT6,1O=R)E\Vg333gbbTWe[[X+GJ-7>,(c=8]OS)5N0@
WbEHW.P0BN_Q;F9W505RH5(>)TFbC>?)8fX8_H4a5J@<XGRZdWaSFJ4V<Ac<fYY[
AgA?O<?:::3U]F,-K,O2Ee3-g8).LFe>E10D0/I+-/U^(KOU\:@Z[4AQ]UXK5^c[
VO>^cCKRT\gB>cTLT8E15CgQDZa+6OJ\Fg6^WLWRNAB(?eX[VEc[(?JG=[,\HdH5
g#WPb+K=)WB[LL^.,^21N949[=CT,-=6B>.IZ0N+>XgMZ6H]2M<J[-G<>F+fg)3,
b-[?Fe;]H&I51K4dX)dfA4,B,&8Bg5/4^8J-:aLRd+3;5\a-?g4PIP[Lc=>3D]Z+
dL8aN&gX&:;/<Z6&1Z/1?NcD6(S4+gW]dM@fAE&P#BH89.]@5A/C[6VT3H]>&DK.
5Z\]E0[3A0X)6EP?e-GAPJ@cXbJ63IM[c>W9Qfe.GDQGK;c&:N]J:J+;MT+0O67L
MY<N(7L5N[/f7@&M^XU<e<.^HG5&V_fa,<S?]0VR@adS\.,D3AXbQ&[N5CZ4[d.<
\3F(TXP7DBM_0NIE;b<BW,&EPR&G-SD<G;a:^Q:1<HSYIaVSD4BC<HG#KKf]#+FF
NC]56?@B2QNOcVV[[NG39S?5[W]/=\CT81CP>K7-80U8G(IKG6_-.OecI#ZX2:M+
V]d\/P7^&K^EOI(0318+)1_:cGf:4fN&d\2U/#MZVFQdD_eX1b4J=0RB#e\?CJ2^
Q;W(1MUe>\;6U-4#N&,8^P&0S;8b:4@Y@NcV_5K85-A8&@W^&>G#K6L+1NT>UXQ[
E>7U01F25Jf+CHE:Ia-.SGcFMbf9/VRVd=Nb1]H]N\d3e<Z>UNb_.X.cJ@R=UEQc
E+35<0PWdNN&0RW+cfSc_O@50M#UcFXT5R;G42FdWH)PJf-7QCeH9_&&Zg5SSFNM
OUUM7U/=T32[D83P4f:1aORQJ.@]/:ATeGL6fO)?Y9HQcI+NH?O]3K:gIb1]V@3;
K-RFLf>)b(7.0ADB>T4YQQLZ9G1^gTUb:K(E#g:J3:J4.a/MJU;+(;2Q8GI2N=)H
A[L:515D(>>B-Ve-113?/<fGKA=.2?BAJ<GXL#32+bfH[0F8bONKQL\gWbJOe8;#
BO<A\T2[?46&1D3-IHN5L]E1;3Gf>)BL/8HY=BK)gW9A#_?[CG7W0ebG)4Ngc038
)BbAT5^Z[7+b#QHdFKNUU009?-Z&(049LU0U.S@[HW>?CX^VYDQ+bKNg7E_MA)I2
aPg<X:OgMNfDGe079XJ1QY4N?TIBGe4<P:T&BSJRBPWZMNb_6-_K=W6QAIBb8^.H
HXG_FT/=.CAcQW6.]/J6.3R.=b1XYZBXWDQIXA:<U_R#][J,LN=+:,8f=L=Y[F,K
0fOUC90Q\ZW9Z(K=M,?VQC\O>>&M:VCK-J+/9@(DcGX_[.Q=9)R(4REPIEV3.<7:
RREM:3JXeOWa/N9[8f67^(Q<>fD_.bMT30SIRP_bVM@BJ+>bH0RALXf_2(>9.^Ng
Ac-a4GegcQR]WKa]X>/?20@7M).]DE#Y#Na5KD.9V8f-H:D3D2?>3Mf)4J:ecM]V
9@/L6>A?K12N&)46S.H#dfOUgd3/<H&@[[=].M_4Aa)-IMX@<T7E7:5),)P<TCF1
KCD,ILA4_G8[ERU(3XLb(MT:9&L+SBB#MKcC3,b7BdVe=&dLJIb4d7=W,c5=HUg_
O;3CTGV6c[M,#]aC1^SQCL-MK^Ld@:#J&NE9#T8;6Cg5)0D]QRLY/8OMbQY?V<b1
H^)H/0?1Z9-@YH.UMXaC@1KYNX:K=_S#3U;Gd:M<ZJM>(</5GM:B1cY(9f:E]##H
7B0AaV&2S\LQRPF[OL/?F\Q&QZQ[39+NaY^BO(G[=,9eL.M0#9bRUcF+T#8Kg+WC
088Ec7bY/DJVPXX33f_-9KP?&^)L?K=M@EX1VH\[YKOBBP-HWWb4_P)4N4UOSg>/
H.?T#KT#Nd?L.<).0(L2(R=C&.6@#KJ99NFU(-Y/-XO52Z?YIJ9(KdYS)#&DV7=U
#)fWB89;Y/8.27N72H4>.Q7FLWA&B@IRP#Kg6>XP&[4+B9WVL#7C7G2B9^TPJ(U<
<TA^e3+QH2E+SXV_Ue\H8--YA&3NSREB[X]7\2DHQA04/H^].g+RAL\Z2\G<Lg2[
GAOKHIKMA2#-U,EVQ6_?M0&XN8#E5\fKG;Jd^[#@JHQD2,:N-JR/PC.@;>2-RN^L
4BNbSDN]DP.^543??Z2NEUcTcE;F?f,RAO3B@^_([)-T36XaM)#[OfE)=g1S>]6)
G>LI9de[;d1EJ<T,^^3E2]?56E]f\3[c@PTH<&(3J>FC)JQ0[@FLCWbfW[Z7+#=#
H+T^]SC.c:J17XD/G1TZ(1JbAIc7b@#0eeVE-&W8XB@.?F1MIJ<@&(=X>5VX)F&S
HS6g478PIQCL8-86@/0TVRM,>]=A+HKF[GDKNARHL25IOC9be>W/=LEa-<J8>,=d
cP8:B\C^7dX)@>[IBAZOZSZ[7Z98SR+ddNQ30[)R;RKeY0b_V?3:G1^4b)C_QS-0
)R_9>]JV3]>Y=N.#\N9,7\[,#Z6=:I5.<G1.KM5X\&YL-NX_HQYcaZ1cMI2LRAXU
>@^)^PC+>)-K&[E/aQ&^&79I:O?Z@ebb?KJ2]6NeS.EC>&YW>#<BL1+U0b26a]P5
O8D<G-bgOYbe)^3C[W70M#J=<M+8=Zea^Id0=;bB+39aC\B^BR744IWI@6GU>??>
5+TMP#O3?7>4PUc59=;)T63)bBK;,++8Te+[3U96S8#4GAKFLW9;)<FA8a#]KaJ6
1K<b\L>;(#(XQB:g[65(H32g-1O.:DJL1+&g?E_W1ZeQM/E(:V;45gIbGE_BKf?D
a_Pe3R9L(;2HL9gbT/MHD3)>TQ<&a<(O5@Id<ZAd0eSOQc8SMSGQ#I>NW:?79S8C
3.X)_Pg0Adf[7fT)><Y(WLd.ID;X2_MBRHM0^0ZI]7H]XQ6W<g))CI+]PA<&Z&c1
(1.CR\d)\-#(G3<^c>V:NVMKU>aecD0Q<8.SCBT&LG.dAgTeR-gE_^TL:\Vc_[CB
Wdb5P,K;]0)Kf)@e?gZ1A8H6U5,#P&^H#LBZ\c@C&VMHFGYDKL2M4CTO0M[=IUB-
\?NYSZ36XW4+R_bcDY)Oe5CD1>H<02>B^Y1PNc;d9#D^FAJ;cEF9Z;[?c/-NW-Z,
-M5HJAE;)eOFNMe-R\KKW3J,2bNNT7JdHJ;R^:&^B3?<2Ub.BQ[D0-?F7-)]Lae-
[);CN:7]Q?AZ,VVK()Ygg\C5=gKYf;P#YY]/P1\0UL8)c(J=\A[GV2I587S?1+<&
Z.VN+Q^L_1I2eVG,SV4KDaR)_)2bI9LMRO-W;DAPE0B4\2(I7/3?_c;cD)SSedR<
:@I37K+M,(.UWg1Ie+9.b/?#6Y80[L&a=5fEQ@EZ4X/NG4A-L<RE:g2U0OCWa@YI
Tb^378R\BEM]4#b+e>[;7c:X?-5P)]?:.5a#OR=__]>e1LI)6fWK?gT2e.^>B3?Z
;>MDe_6CgJR./K(#db/\N&^@e4/S0[)A8FQSe?[K/^H+)6EI?g,AZ/@=VA2LJOMN
-I<>JVA][a.APc.e3+,X@06]<G?P)6gJZ^ID)fF1g.28GU:#5+0-(a#QfR#GPQHG
5H.<UQ6Fa?B@aRYS9&2B+;G+@OE^K8/#,]4>fNYLZTPD:>#\&W=6HCMVI95g[Z&#
&N)Q]HeA2g,\25@OX&4YF,gM2O_4f-BbW6NJ=EE((MQ15ZA.,d5B)f&,.4@SZ+YO
5aY;EV[^2?A>>J^5cM642>D=9T094WL/D]()Y6NfW0Sf7Za=A>a3GA+@Kg1^G6H8
g^2)W&&4@C_RTQR@(PH/OIK#NM0V[1aC20>86B3Oa20^UcbVQLBbZD#d.4cec89W
:_[U)c2Ec=]&gCASgU5;(T\d,<=PJZHD?OMdIL.d<a=]G_5#ffZ<3=TVJJffRG^E
R>fLAAKN0OG\G=-[M;4#3E_C&R)^.<(W<adP@W_J:G(_ee(_5EG^&(O]HR_>B/D^
:PV1GQ^(IS,WOIYPJRg>)#+NU@6RI_PIE1QS,&4aS7_V7C05V#P[)7?VS/Z>K8JR
UOR\eP8[F[K.TH26+Q1X4fO[2Lc4+I@QM-fcQAE3=?[15c@@1JR@\6V43K^;?]e4
FA[3N/&.I@]V-@<03F3f=a0S\[<[#MA,a:)W[M,fL3UHL2PAUPME<&#R<S\+3DDE
A:O_IDKcQN9/Oe]//._H2P\#Z8/@S_7:Q@),L6B4@&YW&-J;S\;#c_-?;>>4>e.Z
.J6N>,EWCS9-U7)f<_9_=;8H@1CRB31NXbX\/bfDb(W3)(^@:c9EAA-/ggYCG?\-
5/HWM9E96.X60783I03I8EHKNI]aPNc_J@)+IdZQ>dXe._Z3G]4BcS^.T3Y,8bD=
g56=G(_+U,-M^WT3CNdM#=[)Fg>M1W27GbE<6QD?)K,=:N2fcTK=&(P7>CEMa=OQ
9]X/FP>1RcHaEH+#.]f5CTUAN45gA6LY\ef@C^Z9Ed2[>2.^J&B3b2DC?Pb)3Ef_
N2IX5GDO^<4TLCB;A_C-BN/,,A0bB:JCbO4.-<>b&B5T5/cMUB=5X52AQ[TfZcd&
MMHQBV33/D&<:K7>=)U[aDOI3JeGH59^=0U9+01PX#(N,\9^(MF#0B&&@dC#L&(U
TA./cYb,V4)-F0(I2b2[:Z\/QgY-D__1<QaO?Ze^(UfC53\U3[0/E=-G@f1MgJ8@
&-T+^[V8Q]aFMB7Va?eHVc(G4c_5[9)(:3;WdcDS6Z,=/J?+Qa>A6YT59e@8PVVa
\I=6I8=[_5[M8>,+\FR=T\EP^6M&[fE_?bFP#6Of9aPF\--]20e&H)Xb;gQ,J7B/
RaZ3H/4)Sf:EV4#1SCd8B&J7Q=g2[-5b0>S;XV)2Te/SXcMcBdZLDPLHZ.7AYQ_#
efPOJU_g)ONWcK8/Oc-].PGLNWFWKZ:aaKY[4K#BE0=I\J4_J[7IUPe3IX3C3^-Q
NX((7G^KVe?N_7dOJI3]S3NPU-^P48W?fS3:=79=:V55dSgFVZ)ABY;K_ed/<OBL
77g,]V5c?\:S1@6@2KJ4a/dVE=a&98WFO/)S_KC\<+N9<^H5(FPMc,Eb:_/UQ1>R
P;85#Md)]J:S@+L9=VQV3^R=59TC[,2F]<6UEKJ&L:]9ILB@^S@4CP2X)a2-.?KW
BNFA+7&f.FbF-_Pc3?J.K3I10WJ5#Ie?0#7.I1-:L#7&]=2E6TbI5.:U\,c.;(4>
c4)L43Z&dCcE5Rb0g+dF5=dWBEB9<>gV20WcbN^(DDfEg=^gYICR?C<5UABb&>3Y
.J>VTaA5S]>:aW]1b7368;9+\K,Q]?S_2UMMd-5VSNYL,6#V#.:d.\+\O5[6daP,
K(d[@MS1/Z7O9cTN5gKU+_7/J4dK<bZW.QSddZ\(W-RC=R\5-85GTQ#^bK.ET8)1
b\2852NT]99S;EOT4YS6_/S]+[Q\9(M?adZL/?:9NR[PJU5@A5W>HeZA:M=<,.8A
KA1Q7:[PEfG.QBFHF<EZ[T2c^gE&Z:L4_CH=PE7Gc4BZ<=<AS@e:/9[:RX>0#@aa
:&J;;^NKA-Y17E#6(@2N;gE+)PMP;(7.8NIcIT:6V\2:E;PQM=@V\UP-E6FIW2>:
6)U[,JWET:TAJ1)fD6FL63=1W2\(4VN3SZDWSE;aC41.I7JP=GT^)5D/,I0VFY:V
#D:C5-^K5e2+&fb.,TG(_#T6:Mb@^9W+F+U;^;FI0T#fT;5ZMGJ<@\LK73,OPJ1T
[8Q;MMR#R.M8MX^DLVK-d&A&3/8eSX,=[fCaBPWP_LS-#Id:8::)F13RJZ:<Jf2:
CI^&c\)01\LW9)d06C9,T^GcJ^d;>P;&EGY:BfSZ//ZX(a=Q0)K[\:[.F,)Q\?A2
8T>ZE>,g;gM\N:MFE@af.:+QD:]A\L\fJ&:@Kf[3C<&HB?LO700@2>PA]<6e[1/_
@84+5I,eg_Rc\^)e4b<UUO_FZf)OA[7)D^.NWPK.MI<.KSGYBPMeDZ^H\NCa\^RL
e^JH7SBe+MJCCg<GFB##ERc@T[B]f?]Dd13+PJ@E&-+.SPW2R?c-AgJ5?#IS#;+]
fJPa=&[=gLO^H;88I/XQ28/D?(N.2S+AL>U1gQ<1OXTBe=HQ#:B<W8&+8AOL<N&8
D;,LX^DZB-M@WCfUb:4B=26,D2?BbM,1_YW4^8c7R9Y&(4#Ac@ZG8=:GOS&A+XTF
YLd-2/I>SG2TZ9921d[1b&./3c&e1AG[fEe)64b1/bJ)4&ALcTUWUQBcR2C]7E]F
F(W\IHf&<UJPJ734feHI];^QN(Z/)JTF6R9,_OB[T0G^2:=WI(@bLSFd7VRXD0G3
;eC8g0)d3DF5b\[EfMFXOQ52XdN)1IXQG5DfG?>HRI&/0QTIR0Zd38W\ZCTQ(e22
SVHN_0TEJRcbJ8bJE;1Ua0S1JKE2UZZS8>7a,@EF:2KZ.:KEADd[8LW+S:Q?IOVg
fdAQdF/4gRR=O<N+M895_6+4aE:[R60MD^YR-#2=@BeSg26466Bc_LC\WQT,/?72
cG(DPJ.QG@aWNE#aA7Qb9,\J\IH=2OV>0XQ,9S6C4@U7N3GWPF\\Y04+>[<:XdeP
AOb1O4,K2MA@<L]Tcf[b31)BTL_@U-\B&09UeQPC>P.E2D-RM&A>SPW^4Tf__,;g
(;1P:_SPBgQ3e9@)2;2H3IW^Y>BJBW3QB[3>QWfV4RL_dL7bT5D)4[2@XW&5M0K<
3^F\GQd,c7B\OY[,DQ63AZb=,4]ZYA<F^2JPX:Yg^ea;^0e?5:TfPG=1G=8E:]9b
Le;GP8EcF@CPNd9C&G8Gg,HE2Qd/X^9DLJbWR7SY9U-Fd-^0E>.ee_6_XWDU]>SK
20aYeU2<7W3WLB9-#d7-IPE\-Fg8&_:PN1FM1NV]aHFac>/6B:.Bd::7>,>^DO^1
2FeQBRMKf/2dZ:)@UA9[Z(dTC4L>7DU_K;RU-J-Z<1XX:;P0eXD.e2EcX;S:+(FT
6&gQ1H0JF\?#g=cJVYKSZ-EUM;.4ST<QM=>&[^dc3>Wcd.=)[[c#1(NP]>5H6>RC
TfK;_Y<6+HaZ@:KY+>5)[U2<Af<JXIL#A2EPcA&7_2@#MST.FgDd?J[Z10B@d35]
\-(RKRZ=#C#W7S=^.UJ(<[R3H.c#GaWC.LTG_]DDO(=2^A(/A^,9,,#H\Zf6RdOg
&VQ7(]-Xd2RN-J28.71#Y(3\#2ZUM([e:/dW0^;(@7R_dGB\U:22L<V_5Be).OU9
DG:V9C3HR+7BJ2GB?H_ZV/J5/N.T#fBKM_J#eFfVPO:2UR#2NWV#LBE#=_VR<KZP
,F>D:F3ZQMXZIQEEDRe15OX1Vb,Xf@=Q9TD9387UU>=>/?G6D2&)Z3^ECB]-^>aV
T1f9<Y^;2PS#QM5deGAIN,ECFO]DA=XC&]BD,C6_B+HUfF5+&FM_@&+V2O89G;eL
&KC^N]@_a[<V.#4&RWa)A\?E=\bI8;YXK6G&EYeQ,AAW4fIeU&H##PH@I/Q\[3Q:
c\g@a]YZ9C(RO5L&5&C973/[KYX4cIC;I1)_=G_BOR3>&UP7P^0f&L]Y948+fZLS
J)e=]EA5<KAXSACX<Q24U[(cU>?;O-Q:EQcfWKdKOV,1K<TR9>VH#e1NK6;[@S<K
_WNPMaQb?)9U1b[Q&I7X>Nd2Z,Xe>877CfcgS.,<gIeI(>1Z8NKADVBPKKDR)=VM
VdB#M5HG9:)AP,_G8YLD_]-1a0W0[Wg2cEQJ_#7XZSJT,CR?]#@<Ge:TP7@FKX0R
\2QI(:d/D0\ZdcYK6N)fJA#,>]QH0bfIL.JBX2NOI5X[Q?ZbO>Oa_ITWI-1d5@/W
5G5D+D]SK#G)^^Y:D8N3@(a(#g^>Bd&A8YK58HKOVfJ@HHB>O4HdP]eYNb>C4;b1
gF8N<@Yd78PL,Z+C8+F^.eJ^]_6_(aWFBC,3C^ZcNH)<c2R^ZU?ScIG^CC;=-7<K
S:@HP(AHa:,0[9b==J@=TN>_STcdd^d/8.Y)P\0D[O925I2g>f,HNfT1L>^L3M.3
9<WV<.g49g[YM9;@g>\[_7f:\?OGEg:^4a-/2g<8cGWPT=XWf^5Z;KgB:gb\E&/F
T-WG/9^#XFI)#WGF_R=IVbHM75GJB[Q]8b4DU_6DaH.C5Q:Z/)US,Zc4]T>:ECCd
Ng^C3=3?B6V@].6H6T1[dS).)>S29:GY;)e0D,XDNbQ9Z<8/:2@gcOc8Fg)cUeg?
CG9IG0ZW;a[XF]DYaQEA438dc30[.E:4-1H79;?(9O&^CAA(<<P9)T]>7Z:.dF<T
46dBUAfbdN&E,.^(]&);BM>acY83_JQ\V;KGFQ+2@<=819.OfKI0d7<Q=GG@MM91
H/_G7DROY\JHgY0@^NMNTMTg[>YVDW>Zfg&.#J\3H8fZM>=&4bQe#SQY@S;f-4&/
>V+33E/X:(WF-20)K3&JBV7fX,6P^]gK>8]9a61D:?G>QaHC-GP1(IS812-)ZH8#
?(0Pg3L9.gZY(OT0(TD<_2[-7JW0BagNEXT,>X^_:V\@#+#^:HH3:?BX;c(DcG04
DfGD[2:RHLEFd8CVQbDPg18165.fcb?#/?GP,?N0BKf.;(,S@ZLT(1:5GeS.7[g#
M3[UXc1E<H)?>A^b[KPKW#=dZ?Hf;[0BU.#1GL/;(Q,I/HR(M5bM=P,)V(;BCG]c
X5H[/bTc3ILJ./FgEY=A-fRaF6b97F<)T1Y&fA4G_H;YY>d>Zc1:NG:243E<4:3&
L:1^SZ3=WB7C1ER(6gc?+]_d3dK^)A.CIV]8A.5=Lc>&\GK@->15\<7I+;f2,L:A
;f?T&6BO6/G0-Yac7^-:a^FVQ#g@aHGIR_-T=@(TL=M(/NYI3HK[URSRH@8^=L?]
e^BRPE1=bd\B^=^.2AbVcMWD)Y>NFMQ5fBX(RQ^<<TRN9Mgf8X<L\ZP41I<C[5EC
2#J^f\)>P.c37X>)X<dD/c?:)Q/97TO[CHGg-Gf_80.P80<U@1\\H?KHHS?&#&BS
IYE-=/cE]JBaBW_FP,;PHYPELC>DVAHV96;^5KLP9dVN2:8L.G--K)3:8.WC[-O-
HLb=/I5ECc+4XIf]0K#.[I8GR&=M\^UQP>C,J[P)F04XSX\+c^^/QK+J^B6Ue^@R
<U_24Q,0Y;@X^=T7fNcE157_-7\DL2Wfb<+Y:<(/;MHW)g[;1N)R8KK850AP<CB9
B]B[AKgSQKMEKP??2;PJcg_74\#F_KJF;/]V#OO#L-W.NY2@OS>,G_PPBZ,X8>RK
/ET;b5?cS_;A:-]R]A&->bN?(UH366@HF7);(BGKce\(B\6W#SKT:.62?gJc3dTR
b&5\++[Y>Z4_N61=;2?8I,&L<7O68XJ:.#:NKKXICI.F,]S5BO=QK()afYSYZdGJ
7->2-[JI.GN^X3DW?2/],V,?:9WfXSI/RLcPHLP/QV4;9N^ZW1RB+YR@W+M9TIXa
]6FgX</\1VfAcZ+@,D7HU51=DIW@<WQ7YDXY^]?))@Zb/=CJ;Be0.3#WgeT=[@HH
[1IWd/W,c^VADYaC:0U2V1[IB,&@[9abBK0#@I(fF-A[ed,[/)T=Q>29]]cbT.)P
9OV^5C-CA6^H,a89V:G;Qbbc9Y+^T1fY;56OL<-OP:H.-g1]aOBE<LAX+&Z[6;XW
73g05QI_+B^J6F55),@[[RW9S:6XCS?G7OGTEM6gV]/V/0>\_J&9TaBG-E-aT6J[
G]4OP1,AN5Y1P(UU7c7<&9YaF#:]\4NBPF_FJ+f,Me2#<7[_M(<^R_\I:)-VV6AF
<#:^ETd2@]1E>SP-&>10C1K->1;:VI48E\T,)b95bQBQROfWS6WdKfM.D[;+3e.9
2+4=L7adI.PGA/aXL,(=LZL62Q9HAV_6(HFWRY(:/W-E:3+#4F[/PEEd,:LM_7Xb
T5?\0Y&_U-(PP(&U,K,[aOYH;U+&gCN/Q/+OR^CcdbG,^-1+-f_(][eN4fcb(@/.
1Tf7c#&]Td9/J4FFIPWM]P>d1@-=2&6V^.?;QB=/dgKXK,DJBRFSX1^,]W)Lf+<N
XCJ@NWfUVK\Y^Je8@_AcCaffdTEINfdSfET_d8P@U9R_BC_;A@A5Sa3T54YJacK&
8+DPY\IH33Q.WYff>G:AN[?P?_QF>K:a\HQO@OMH;H4/JA2Z\fb\6\NK7eTYMA/@
XCC><80VYCXZf9]RHQ&NI<4O?/J+C,UF<?YIQa57[;>^9GBGUcVN:]VLJTT8\eWF
>];[FM=Hd[&LWG?I>?P\\D)&=P<5I4-Z&(Q@BDT@O.PG=)76@egY9cVadWC18&2O
g3T])CM&VGLe/>\R[];UC(2?<L6V(_\JSOVC_dT-#\a:F+;gYGTUD5/0]]7_W)S(
?=F@bT.=OM1#W7M@&2])POf(@R-WC4(W<PA6e1c,YgS@eK3:#(>WfI:-&48QE_^V
=6T0/)A6G.UL7)+_JZf4fJ)dVH3D@U,\/d7e:,=7?AA\;(d)\T.AQ)./2LT+NJB9
]4^?XA,+:10+Tb61R#KgM>3GK5/E[C5R[AJg:8+R\[R9(5<dC8@c,2/TeE3>L?P^
MPW2GSIC1W^bC>C]U\MX4gN:IcfF)__4:>7ND.>1SE12B,cMHE_BWB#TE@?e6IF+
1]52WWI[M@U@;EZIJ8,#fD7OHR_>0-HGaBXR0P;Vg/VQa5\9b2ZG-S=__2f?G+KP
[M--^a0HS?2C56N5U0,cXA]Ye#F#3HGBa5YR@+W4+DH0d(]DQ)W\F@fW4ZO,:=+S
TQI<//Q[EN>?DJae9)3T[(ZRe?b+9XV3#+4^I[QM.NZIM@Ad?[1[1+@Y@SXaP-,M
ZC-SF&Ob[TT0,b4^3/5UV?EBFI3I7Q.R5^b-6-B=(D1OMf6<d/=8Bc<T:6NUIN0L
e_4>Z6P.Y2IAUaQ93eYV]./PGSFPVO>+e17\F_<0XW76/L/AM+QfT?]:#<25:-AM
ZH.8RYGMV8bUXd#API+J(a2SRUIAK1@.L_LDS@XFB.4YGIQcRf.a^T]?Y1>D-d(O
NXM\e4<)/TH=LG.JK@>Q8]2S6$
`endprotected
endmodule
// ##############################################################
//   You can modify by your own
//   You can modify by your own
//   You can modify by your own
// ##############################################################

module CHIP(
    // input signals
    clk,
    rst_n,
    in_valid, 
    in_valid2,
    
    image,
    template,
    image_size,
	action,
	
    // output signals
    out_valid,
    out_value
);


input            clk, rst_n, in_valid, in_valid2;
input     [7:0]  image;
input     [7:0]  template;
input     [1:0]  image_size;
input     [2:0]  action;

output           out_valid;
output           out_value;

//==================================================================
// reg & wire
//==================================================================
wire             C_clk;
wire             C_rst_n;
wire             C_in_valid;
wire             C_in_valid2;

wire     [7:0]   C_image;
wire     [7:0]   C_template;
wire     [1:0]   C_image_size;
wire     [2:0]   C_action;

wire             C_out_valid;
wire             C_out_value;

//==================================================================
// CORE
//==================================================================
TMIP CORE(
	// input signals
    .clk(C_clk),
    .rst_n(C_rst_n),
    .in_valid(C_in_valid), 
    .in_valid2(C_in_valid2),
    
    .image(C_image),
    .template(C_template),
    .image_size(C_image_size),
	.action(C_action),
	
    // output signals
    .out_valid(C_out_valid),
    .out_value(C_out_value)
);

//==================================================================
// INPUT PAD
// Syntax: XMD PAD_NAME ( .O(CORE_PORT_NAME), .I(CHIP_PORT_NAME), .PU(1'b0), .PD(1'b0), .SMT(1'b0));
//     Ex: XMD    I_CLK ( .O(C_clk),          .I(clk),            .PU(1'b0), .PD(1'b0), .SMT(1'b0));
//==================================================================
// You need to finish this part
XMD I_CLK           ( .O(C_clk),                .I(clk),                .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_RST_N         ( .O(C_rst_n),              .I(rst_n),              .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IN_VALID      ( .O(C_in_valid),           .I(in_valid),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IN_VALID2     ( .O(C_in_valid2),          .I(in_valid2),          .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE_0       ( .O(C_image[0]),           .I(image[0]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE_1       ( .O(C_image[1]),           .I(image[1]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE_2       ( .O(C_image[2]),           .I(image[2]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE_3       ( .O(C_image[3]),           .I(image[3]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE_4       ( .O(C_image[4]),           .I(image[4]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE_5       ( .O(C_image[5]),           .I(image[5]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE_6       ( .O(C_image[6]),           .I(image[6]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE_7       ( .O(C_image[7]),           .I(image[7]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_TEMPLATE_0    ( .O(C_template[0]),        .I(template[0]),        .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_TEMPLATE_1    ( .O(C_template[1]),        .I(template[1]),        .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_TEMPLATE_2    ( .O(C_template[2]),        .I(template[2]),        .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_TEMPLATE_3    ( .O(C_template[3]),        .I(template[3]),        .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_TEMPLATE_4    ( .O(C_template[4]),        .I(template[4]),        .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_TEMPLATE_5    ( .O(C_template[5]),        .I(template[5]),        .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_TEMPLATE_6    ( .O(C_template[6]),        .I(template[6]),        .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_TEMPLATE_7    ( .O(C_template[7]),        .I(template[7]),        .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE_SIZE_0  ( .O(C_image_size[0]),      .I(image_size[0]),      .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE_SIZE_1  ( .O(C_image_size[1]),      .I(image_size[1]),      .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_ACTION_0      ( .O(C_action[0]),          .I(action[0]),          .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_ACTION_1      ( .O(C_action[1]),          .I(action[1]),          .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_ACTION_2      ( .O(C_action[2]),          .I(action[2]),          .PU(1'b0), .PD(1'b0), .SMT(1'b0));


//==================================================================
// OUTPUT PAD
// Syntax: YA2GSD PAD_NAME (.I(CORE_PIN_NAME), .O(PAD_PIN_NAME), .E(1'b1), .E2(1'b1), .E4(1'b1), .E8(1'b0), .SR(1'b0));
//     Ex: YA2GSD  O_VALID (.I(C_out_valid),   .O(out_valid),    .E(1'b1), .E2(1'b1), .E4(1'b1), .E8(1'b0), .SR(1'b0));
//==================================================================
// You need to finish this part
YA2GSD O_VALID    ( .I(C_out_valid),    .O(out_valid),    .E(1'b1), .E2(1'b1), .E4(1'b1), .E8(1'b0), .SR(1'b0));
YA2GSD O_VALUE    ( .I(C_out_value),    .O(out_value),    .E(1'b1), .E2(1'b1), .E4(1'b1), .E8(1'b0), .SR(1'b0));


//==================================================================
// I/O power 3.3V pads x? (DVDD + DGND)
// Syntax: VCC3IOD/GNDIOD PAD_NAME ();
//    Ex1: VCC3IOD        VDDP0 ();
//    Ex2: GNDIOD         GNDP0 ();
//==================================================================
// You need to finish this part
// One power pad can provide power for 3~4 Output Pads or 6~8 Input Pads
// We have 25 Input Pads and 2 Output Pads
// So, we need about 4 power pads
VCC3IOD VDDP0 ();
VCC3IOD VDDP1 ();
VCC3IOD VDDP2 ();
VCC3IOD VDDP3 ();
GNDIOD  GNDP0 ();
GNDIOD  GNDP1 ();
GNDIOD  GNDP2 ();
GNDIOD  GNDP3 ();


//==================================================================
// Core power 1.8V pads x? (VDD + GND)
// Syntax: VCCKD/GNDKD PAD_NAME ();
//    Ex1: VCCKD       VDDC0 ();
//    Ex2: GNDKD       GNDC0 ();
//==================================================================
// You need to finish this part
// One core power pad can provide 40~50 mA current
// That is, 50mA * 1.8V = 90mW
// From power report, the total power is 24.0552 mW
// So, we need about 1 core power pad, but choose 2 for safety
VCCKD VDDC0 ();
VCCKD VDDC1 ();
GNDKD GNDC0 ();
GNDKD GNDC1 ();


endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Ultra(TM) in wire load mode
// Version   : T-2022.03
// Date      : Fri Nov 29 19:43:20 2024
/////////////////////////////////////////////////////////////


module TMIP ( clk, rst_n, in_valid, in_valid2, image, template, image_size, 
        action, out_valid, out_value );
  input [7:0] image;
  input [7:0] template;
  input [1:0] image_size;
  input [2:0] action;
  input clk, rst_n, in_valid, in_valid2;
  output out_valid, out_value;
  wire   mem_we_a, mem_cs_a, mem_we_a_reg, N442, last_in_valid2, action_done,
         out_valid_a1, last_in_valid, last_in_valid_d1, action_5_flag, N7421,
         N7422, N7502, N7503, N7504, N7505, N7766, N7767, N7768, N7769, N7770,
         N7771, N7772, N7773, N7774, N7775, N7776, N7777, N7778, N7779, N7780,
         N7781, N7782, N7783, N7784, N7785, out_value_a1, C551_DATA2_0,
         C551_DATA2_1, C551_DATA2_2, C551_DATA2_3, C551_DATA2_4, C551_DATA2_5,
         C551_DATA2_6, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, net76341,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         C1_Z_6, C1_Z_5, C1_Z_4, C1_Z_3, C1_Z_2, C1_Z_1, C1_Z_0,
         DP_OP_989J1_126_3015_n7, DP_OP_989J1_126_3015_n6,
         DP_OP_989J1_126_3015_n5, DP_OP_989J1_126_3015_n4,
         DP_OP_989J1_126_3015_n3, DP_OP_989J1_126_3015_n2,
         DP_OP_989J1_126_3015_n1, intadd_204_CI, intadd_206_CI, intadd_1_CI,
         intadd_2_A_0_, intadd_4_CI, intadd_5_B_0_, intadd_5_CI, intadd_8_B_0_,
         intadd_8_CI, intadd_11_B_0_, intadd_11_CI, intadd_13_CI,
         intadd_14_B_0_, intadd_14_CI, intadd_16_B_0_, intadd_16_CI,
         intadd_19_B_0_, intadd_22_CI, intadd_25_A_0_, intadd_25_B_0_,
         intadd_28_A_0_, intadd_32_CI, intadd_36_CI, intadd_39_B_0_,
         intadd_42_CI, intadd_44_CI, intadd_45_CI, intadd_47_CI, intadd_48_CI,
         intadd_50_CI, intadd_55_CI, intadd_57_CI, intadd_59_CI, intadd_60_CI,
         intadd_62_B_0_, intadd_65_CI, intadd_66_CI, intadd_68_CI,
         intadd_69_CI, intadd_71_CI, intadd_72_B_0_, intadd_72_CI,
         intadd_77_CI, intadd_82_CI, intadd_83_CI, intadd_85_B_1_,
         intadd_86_B_1_, intadd_86_CI, intadd_88_CI, intadd_89_B_1_,
         intadd_89_CI, intadd_94_CI, intadd_96_B_1_, intadd_96_CI,
         intadd_97_B_1_, intadd_97_CI, intadd_98_CI, intadd_99_CI,
         intadd_101_CI, intadd_103_CI, intadd_105_CI, intadd_106_CI,
         intadd_108_CI, intadd_109_CI, intadd_111_CI, intadd_112_CI,
         intadd_115_CI, intadd_117_CI, intadd_119_CI, intadd_120_B_1_,
         intadd_120_CI, intadd_122_CI, intadd_123_CI, intadd_125_CI,
         intadd_129_CI, intadd_130_A_0_, intadd_130_B_0_, intadd_132_B_1_,
         intadd_134_CI, intadd_137_A_0_, intadd_137_B_0_, intadd_140_CI,
         intadd_142_CI, intadd_145_CI, intadd_147_CI, intadd_148_CI,
         intadd_150_CI, intadd_151_CI, intadd_153_CI, intadd_156_CI,
         intadd_158_CI, intadd_159_B_1_, intadd_159_CI, intadd_162_CI,
         intadd_169_CI, intadd_171_B_0_, intadd_186_A_0_, intadd_188_A_0_,
         intadd_188_B_0_, intadd_189_A_0_, intadd_189_B_0_, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
         n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
         n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
         n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
         n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
         n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
         n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
         n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
         n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507,
         n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
         n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
         n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
         n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
         n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
         n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
         n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
         n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
         n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
         n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
         n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
         n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603,
         n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
         n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
         n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
         n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
         n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643,
         n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651,
         n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
         n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
         n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675,
         n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683,
         n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691,
         n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699,
         n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
         n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715,
         n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723,
         n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
         n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
         n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747,
         n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755,
         n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
         n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771,
         n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
         n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
         n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795,
         n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
         n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
         n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819,
         n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827,
         n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
         n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843,
         n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
         n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859,
         n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867,
         n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
         n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
         n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891,
         n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899,
         n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
         n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915,
         n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
         n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931,
         n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939,
         n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947,
         n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
         n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963,
         n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971,
         n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
         n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987,
         n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
         n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003,
         n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011,
         n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019,
         n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
         n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035,
         n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043,
         n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
         n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059,
         n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067,
         n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075,
         n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083,
         n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091,
         n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
         n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107,
         n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115,
         n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
         n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131,
         n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139,
         n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147,
         n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155,
         n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163,
         n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
         n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179,
         n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187,
         n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
         n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203,
         n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211,
         n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219,
         n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227,
         n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235,
         n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243,
         n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251,
         n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259,
         n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267,
         n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275,
         n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283,
         n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291,
         n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299,
         n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307,
         n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315,
         n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323,
         n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331,
         n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339,
         n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347,
         n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355,
         n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363,
         n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371,
         n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379,
         n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387,
         n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395,
         n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403,
         n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411,
         n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419,
         n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427,
         n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435,
         n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443,
         n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451,
         n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459,
         n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467,
         n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475,
         n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483,
         n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491,
         n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499,
         n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507,
         n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515,
         n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523,
         n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531,
         n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539,
         n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547,
         n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555,
         n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563,
         n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571,
         n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579,
         n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587,
         n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595,
         n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603,
         n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611,
         n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619,
         n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627,
         n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635,
         n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643,
         n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651,
         n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659,
         n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667,
         n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675,
         n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683,
         n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691,
         n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699,
         n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707,
         n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715,
         n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723,
         n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731,
         n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739,
         n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747,
         n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755,
         n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763,
         n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771,
         n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779,
         n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787,
         n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795,
         n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803,
         n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811,
         n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819,
         n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827,
         n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835,
         n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843,
         n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851,
         n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859,
         n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867,
         n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875,
         n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883,
         n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891,
         n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899,
         n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907,
         n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915,
         n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923,
         n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931,
         n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939,
         n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947,
         n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955,
         n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963,
         n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971,
         n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979,
         n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987,
         n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995,
         n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003,
         n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011,
         n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019,
         n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027,
         n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035,
         n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043,
         n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051,
         n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059,
         n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067,
         n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075,
         n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083,
         n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091,
         n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099,
         n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107,
         n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115,
         n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123,
         n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131,
         n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139,
         n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147,
         n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155,
         n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163,
         n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171,
         n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179,
         n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187,
         n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195,
         n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203,
         n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211,
         n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219,
         n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227,
         n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235,
         n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243,
         n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251,
         n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259,
         n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267,
         n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275,
         n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283,
         n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291,
         n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299,
         n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307,
         n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315,
         n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323,
         n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331,
         n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339,
         n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347,
         n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355,
         n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363,
         n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371,
         n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379,
         n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387,
         n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395,
         n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403,
         n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411,
         n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419,
         n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427,
         n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435,
         n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443,
         n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451,
         n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459,
         n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
         n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475,
         n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483,
         n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491,
         n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499,
         n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507,
         n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515,
         n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523,
         n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531,
         n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539,
         n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547,
         n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555,
         n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563,
         n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571,
         n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579,
         n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587,
         n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595,
         n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603,
         n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611,
         n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619,
         n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627,
         n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635,
         n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643,
         n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651,
         n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659,
         n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667,
         n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675,
         n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683,
         n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691,
         n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699,
         n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707,
         n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715,
         n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723,
         n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731,
         n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739,
         n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747,
         n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755,
         n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763,
         n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771,
         n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779,
         n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787,
         n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795,
         n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803,
         n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811,
         n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819,
         n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827,
         n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835,
         n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843,
         n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851,
         n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859,
         n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867,
         n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
         n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883,
         n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891,
         n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899,
         n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907,
         n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915,
         n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923,
         n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931,
         n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
         n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
         n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955,
         n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963,
         n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
         n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979,
         n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987,
         n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995,
         n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003,
         n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011,
         n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019,
         n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027,
         n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035,
         n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043,
         n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051,
         n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059,
         n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067,
         n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075,
         n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083,
         n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091,
         n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099,
         n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107,
         n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
         n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123,
         n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131,
         n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139,
         n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147,
         n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155,
         n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163,
         n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171,
         n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179,
         n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187,
         n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195,
         n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203,
         n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211,
         n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219,
         n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227,
         n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235,
         n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243,
         n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251,
         n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259,
         n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267,
         n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275,
         n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283,
         n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291,
         n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299,
         n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307,
         n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315,
         n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323,
         n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331,
         n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339,
         n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347,
         n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355,
         n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363,
         n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
         n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379,
         n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387,
         n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395,
         n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403,
         n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411,
         n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419,
         n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427,
         n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435,
         n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443,
         n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451,
         n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459,
         n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467,
         n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475,
         n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483,
         n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491,
         n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499,
         n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507,
         n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515,
         n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523,
         n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531,
         n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539,
         n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547,
         n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555,
         n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563,
         n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571,
         n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579,
         n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587,
         n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595,
         n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603,
         n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611,
         n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619,
         n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627,
         n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635,
         n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643,
         n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651,
         n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659,
         n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667,
         n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675,
         n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683,
         n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691,
         n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699,
         n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707,
         n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715,
         n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723,
         n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731,
         n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739,
         n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747,
         n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755,
         n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763,
         n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771,
         n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779,
         n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787,
         n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795,
         n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803,
         n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811,
         n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819,
         n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827,
         n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835,
         n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843,
         n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851,
         n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859,
         n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867,
         n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875,
         n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883,
         n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891,
         n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899,
         n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907,
         n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915,
         n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923,
         n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931,
         n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939,
         n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947,
         n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955,
         n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963,
         n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971,
         n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979,
         n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987,
         n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995,
         n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003,
         n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011,
         n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019,
         n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027,
         n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035,
         n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043,
         n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051,
         n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059,
         n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067,
         n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075,
         n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083,
         n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091,
         n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099,
         n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107,
         n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115,
         n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123,
         n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131,
         n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139,
         n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147,
         n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155,
         n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163,
         n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171,
         n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179,
         n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187,
         n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195,
         n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203,
         n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211,
         n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219,
         n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227,
         n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235,
         n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243,
         n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251,
         n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259,
         n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267,
         n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275,
         n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283,
         n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291,
         n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299,
         n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307,
         n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315,
         n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323,
         n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331,
         n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339,
         n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347,
         n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355,
         n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363,
         n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371,
         n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
         n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387,
         n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395,
         n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403,
         n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411,
         n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419,
         n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427,
         n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435,
         n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443,
         n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451,
         n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459,
         n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467,
         n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475,
         n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
         n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491,
         n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499,
         n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507,
         n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515,
         n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523,
         n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531,
         n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539,
         n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547,
         n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555,
         n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563,
         n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571,
         n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
         n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587,
         n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595,
         n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603,
         n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611,
         n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619,
         n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627,
         n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635,
         n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643,
         n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651,
         n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659,
         n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667,
         n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675,
         n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683,
         n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
         n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699,
         n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707,
         n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715,
         n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
         n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731,
         n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739,
         n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747,
         n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755,
         n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763,
         n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771,
         n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779,
         n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787,
         n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795,
         n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803,
         n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811,
         n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819,
         n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827,
         n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835,
         n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843,
         n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851,
         n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859,
         n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867,
         n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875,
         n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883,
         n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891,
         n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899,
         n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907,
         n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915,
         n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923,
         n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931,
         n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939,
         n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947,
         n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955,
         n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963,
         n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971,
         n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979,
         n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987,
         n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995,
         n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003,
         n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011,
         n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019,
         n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027,
         n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035,
         n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043,
         n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051,
         n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059,
         n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067,
         n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075,
         n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083,
         n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091,
         n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099,
         n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107,
         n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115,
         n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123,
         n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131,
         n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139,
         n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147,
         n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155,
         n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163,
         n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171,
         n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179,
         n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187,
         n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195,
         n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203,
         n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211,
         n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219,
         n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227,
         n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235,
         n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243,
         n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251,
         n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259,
         n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267,
         n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275,
         n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283,
         n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291,
         n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299,
         n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307,
         n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315,
         n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323,
         n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331,
         n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339,
         n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347,
         n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355,
         n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363,
         n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371,
         n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379,
         n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387,
         n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395,
         n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403,
         n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411,
         n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419,
         n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427,
         n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435,
         n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443,
         n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451,
         n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459,
         n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467,
         n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475,
         n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483,
         n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491,
         n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499,
         n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507,
         n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515,
         n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523,
         n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531,
         n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539,
         n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547,
         n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555,
         n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563,
         n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571,
         n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579,
         n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587,
         n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595,
         n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603,
         n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611,
         n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619,
         n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627,
         n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635,
         n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643,
         n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651,
         n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659,
         n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667,
         n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675,
         n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683,
         n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691,
         n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26699,
         n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707,
         n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715,
         n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723,
         n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731,
         n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739,
         n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747,
         n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755,
         n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763,
         n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771,
         n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779,
         n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787,
         n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795,
         n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803,
         n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811,
         n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819,
         n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827,
         n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835,
         n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843,
         n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851,
         n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859,
         n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867,
         n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875,
         n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883,
         n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891,
         n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899,
         n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907,
         n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915,
         n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923,
         n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931,
         n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939,
         n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947,
         n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955,
         n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963,
         n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971,
         n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979,
         n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987,
         n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995,
         n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003,
         n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011,
         n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019,
         n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027,
         n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035,
         n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043,
         n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051,
         n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059,
         n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067,
         n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075,
         n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083,
         n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091,
         n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099,
         n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107,
         n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115,
         n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123,
         n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131,
         n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139,
         n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147,
         n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155,
         n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163,
         n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171,
         n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179,
         n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187,
         n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195,
         n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203,
         n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211,
         n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219,
         n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227,
         n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235,
         n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243,
         n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251,
         n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259,
         n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267,
         n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275,
         n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283,
         n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291,
         n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299,
         n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307,
         n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315,
         n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323,
         n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331,
         n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339,
         n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347,
         n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355,
         n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363,
         n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371,
         n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379,
         n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387,
         n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395,
         n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403,
         n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411,
         n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419,
         n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427,
         n27428, n27429, n27430, n27431, n27432, n27433, n27434, n27435,
         n27436, n27437, n27438, n27439, n27440, n27441, n27442, n27443,
         n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451,
         n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459,
         n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467,
         n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475,
         n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483,
         n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491,
         n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499,
         n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507,
         n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515,
         n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523,
         n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531,
         n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539,
         n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547,
         n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555,
         n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563,
         n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571,
         n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579,
         n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27587,
         n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595,
         n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603,
         n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611,
         n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619,
         n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627,
         n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635,
         n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643,
         n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651,
         n27652, n27653, n27654, n27655, n27656, n27657, n27658, n27659,
         n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667,
         n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675,
         n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683,
         n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691,
         n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699,
         n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707,
         n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715,
         n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723,
         n27724, n27725, n27726, n27727, n27728, n27729, n27730, n27731,
         n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739,
         n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747,
         n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755,
         n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763,
         n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771,
         n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779,
         n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787,
         n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795,
         n27796, n27797, n27798, n27799, n27800, n27801, n27802, n27803,
         n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811,
         n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819,
         n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827,
         n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835,
         n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843,
         n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851,
         n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859,
         n27860, n27861, n27862, n27863, n27864, n27865, n27866, n27867,
         n27868, n27869, n27870, n27871, n27872, n27873, n27874, n27875,
         n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883,
         n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891,
         n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899,
         n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907,
         n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915,
         n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923,
         n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931,
         n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939,
         n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947,
         n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955,
         n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963,
         n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971,
         n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979,
         n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987,
         n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995,
         n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003,
         n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011,
         n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28019,
         n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027,
         n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035,
         n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043,
         n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051,
         n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059,
         n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067,
         n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075,
         n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083,
         n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091,
         n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099,
         n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107,
         n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115,
         n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123,
         n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131,
         n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139,
         n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147,
         n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155,
         n28156, n28157, n28158, n28159, n28160, n28161, n28162, n28163,
         n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171,
         n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179,
         n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187,
         n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195,
         n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203,
         n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211,
         n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219,
         n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227,
         n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235,
         n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243,
         n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251,
         n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259,
         n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267,
         n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275,
         n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283,
         n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291,
         n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299,
         n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307,
         n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315,
         n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323,
         n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331,
         n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339,
         n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347,
         n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355,
         n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363,
         n28364, n28365, n28366, n28367, n28368, n28369, n28370, n28371,
         n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379,
         n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387,
         n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395,
         n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403,
         n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411,
         n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419,
         n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427,
         n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435,
         n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443,
         n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451,
         n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459,
         n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467,
         n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475,
         n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483,
         n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491,
         n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499,
         n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507,
         n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515,
         n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523,
         n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531,
         n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539,
         n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547,
         n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555,
         n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563,
         n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571,
         n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579,
         n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587,
         n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595,
         n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603,
         n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611,
         n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619,
         n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627,
         n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635,
         n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643,
         n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651,
         n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659,
         n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667,
         n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675,
         n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683,
         n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691,
         n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699,
         n28700, n28701, n28702, n28703, n28704, n28705, n28706, n28707,
         n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715,
         n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723,
         n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731,
         n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739,
         n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747,
         n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755,
         n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763,
         n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771,
         n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779,
         n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787,
         n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795,
         n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803,
         n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811,
         n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819,
         n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827,
         n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835,
         n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843,
         n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28851,
         n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859,
         n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867,
         n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875,
         n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883,
         n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891,
         n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899,
         n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907,
         n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915,
         n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923,
         n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931,
         n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939,
         n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947,
         n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28955,
         n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963,
         n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971,
         n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979,
         n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987,
         n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995,
         n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003,
         n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011,
         n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019,
         n29020, n29021, n29022, n29023, n29024, n29025, n29026, n29027,
         n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035,
         n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043,
         n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051,
         n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059,
         n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067,
         n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075,
         n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083,
         n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091,
         n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099,
         n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107,
         n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115,
         n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123,
         n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131,
         n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139,
         n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147,
         n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155,
         n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163,
         n29164, n29165, n29166, n29167, n29168, n29169, n29170, n29171,
         n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179,
         n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187,
         n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195,
         n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203,
         n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211,
         n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219,
         n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227,
         n29228, n29229, n29230, n29231, n29232, n29233, n29234, n29235,
         n29236, n29237, n29238, n29239, n29240, n29241, n29242, n29243,
         n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251,
         n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259,
         n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267,
         n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275,
         n29276, n29277, n29278, n29279, n29280, n29281, n29282, n29283,
         n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291,
         n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299,
         n29300, n29301, n29302, n29303, n29304, n29305, n29306, n29307,
         n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315,
         n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323,
         n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331,
         n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339,
         n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347,
         n29348, n29349, n29350, n29351, n29352, n29353, n29354, n29355,
         n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363,
         n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371,
         n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379,
         n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387,
         n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395,
         n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403,
         n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411,
         n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419,
         n29420, n29421, n29422, n29423, n29424, n29425, n29426, n29427,
         n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435,
         n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443,
         n29444, n29445, n29446, n29447, n29448, n29449, n29450, n29451,
         n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459,
         n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467,
         n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475,
         n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483,
         n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491,
         n29492, n29493, n29494, n29495, n29496, n29497, n29498, n29499,
         n29500, n29501, n29502, n29503, n29504, n29505, n29506, n29507,
         n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515,
         n29516, n29517, n29518, n29519, n29520, n29521, n29522, n29523,
         n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531,
         n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539,
         n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547,
         n29548, n29549, n29550, n29551, n29552, n29553, n29554, n29555,
         n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563,
         n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571,
         n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579,
         n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587,
         n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595,
         n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603,
         n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611,
         n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619,
         n29620, n29621, n29622, n29623, n29624, n29625, n29626, n29627,
         n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635,
         n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643,
         n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651,
         n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659,
         n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667,
         n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675,
         n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683,
         n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691,
         n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699,
         n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707,
         n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715,
         n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723,
         n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731,
         n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739,
         n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747,
         n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755,
         n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763,
         n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771,
         n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779,
         n29780, n29781, n29782, n29783, n29784, n29785, n29786, n29787,
         n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795,
         n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803,
         n29804, n29805, n29806, n29807, n29808, n29809, n29810, n29811,
         n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29819,
         n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827,
         n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835,
         n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843,
         n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851,
         n29852, n29853, n29854, n29855, n29856, n29857, n29858, n29859,
         n29860, n29861, n29862, n29863, n29864, n29865, n29866, n29867,
         n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875,
         n29876, n29877, n29878, n29879, n29880, n29881, n29882, n29883,
         n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891,
         n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899,
         n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907,
         n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915,
         n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923,
         n29924, n29925, n29926, n29927, n29928, n29929, n29930, n29931,
         n29932, n29933, n29934, n29935, n29936, n29937, n29938, n29939,
         n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947,
         n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955,
         n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963,
         n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971,
         n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979,
         n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987,
         n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995,
         n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003,
         n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011,
         n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019,
         n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30027,
         n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035,
         n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043,
         n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051,
         n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059,
         n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067,
         n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075,
         n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083,
         n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091,
         n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099,
         n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107,
         n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115,
         n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123,
         n30124, n30125, n30126, n30127, n30128, n30129, n30130, n30131,
         n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139,
         n30140, n30141, n30142, n30143, n30144, n30145, n30146, n30147,
         n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155,
         n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163,
         n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171,
         n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179,
         n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187,
         n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195,
         n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203,
         n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211,
         n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219,
         n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227,
         n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235,
         n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243,
         n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251,
         n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259,
         n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267,
         n30268, n30269, n30270, n30271, n30272, n30273, n30274, n30275,
         n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283,
         n30284, n30285, n30286, n30287, n30288, n30289, n30290, n30291,
         n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299,
         n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307,
         n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30315,
         n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323,
         n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331,
         n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339,
         n30340, n30341, n30342, n30343, n30344, n30345, n30346, n30347,
         n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355,
         n30356, n30357, n30358, n30359, n30360, n30361, n30362, n30363,
         n30364, n30365, n30366, n30367, n30368, n30369, n30370, n30371,
         n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379,
         n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387,
         n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395,
         n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403,
         n30404, n30405, n30406, n30407, n30408, n30409, n30410, n30411,
         n30412, n30413, n30414, n30415, n30416, n30417, n30418, n30419,
         n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427,
         n30428, n30429, n30430, n30431, n30432, n30433, n30434, n30435,
         n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443,
         n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451,
         n30452, n30453, n30454, n30455, n30456, n30457, n30458;
  wire   [9:0] mem_addr_a;
  wire   [7:0] mem_data_a_in;
  wire   [7:0] mem_data_a_out;
  wire   [2:0] cs_d1;
  wire   [1:0] image_size_reg_master;
  wire   [3:0] cnt_dyn;
  wire   [1:0] read_layer;
  wire   [8:0] cnt_bdyn;
  wire   [2:0] cs;
  wire   [7:0] gray_scale_0_s;
  wire   [7:0] gray_scale_1_s;
  wire   [7:0] gray_scale_2_s;
  wire   [7:0] template_in_reg;
  wire   [1:0] image_size_in_reg;
  wire   [2:0] action_in_reg;
  wire   [5:0] cnt_20;
  wire   [2:0] action_doing;
  wire   [3:0] cnt_cro_y;
  wire   [3:0] cnt_cro_x;
  wire   [2:0] set_cnt;
  wire   [7:0] cnt;
  wire   [7:0] cnt_n;
  wire   [3:0] cnt_dyn_n;
  wire   [3:0] cnt_dyn_d1;
  wire   [3:0] cnt_dyn_base;
  wire   [1:0] image_size_reg_set;
  wire   [3:0] cnt_bdyn_d1;
  wire   [1:0] cnt_cro_3;
  wire   [1:0] cnt_cro_3b3;
  wire   [5:0] cnt_20_n;
  wire   [71:0] template_reg;
  wire   [23:0] action_reg;
  wire   [7:0] gray_scale_0;
  wire   [9:0] gray_scale_1;
  wire   [7:0] gray_scale_2;
  wire   [9:8] gray_scale_1_n;
  wire   [7:0] gray_scale_2_n;
  wire   [3:0] medfilt_state;
  wire   [2047:0] gray_img;
  wire   [3:0] medfilt_state_d1;
  wire   [3:0] medfilt_cnt2_d1;
  wire   [3:0] medfilt_cnt_d1;
  wire   [7:0] medfilt_out_reg;
  wire   [127:0] mem_data_out_reg_shift_0;
  wire   [127:0] mem_data_out_reg_shift_1;
  wire   [31:0] mem_data_out_reg_shift_2;
  wire   [3:0] medfilt_cnt;
  wire   [3:0] medfilt_cnt2;
  wire   [19:0] cro_mac;
  wire   [19:0] cro_mac_store;

  SUMA180_768X8X1BM2 MEM1024_instance_SUMA180_768X8X1BM2_instance ( .A0(
        mem_addr_a[0]), .A1(mem_addr_a[1]), .A2(mem_addr_a[2]), .A3(
        mem_addr_a[3]), .A4(mem_addr_a[4]), .A5(mem_addr_a[5]), .A6(
        mem_addr_a[6]), .A7(mem_addr_a[7]), .A8(mem_addr_a[8]), .A9(
        mem_addr_a[9]), .CK(clk), .CS(mem_cs_a), .DI0(mem_data_a_in[0]), .DI1(
        mem_data_a_in[1]), .DI2(mem_data_a_in[2]), .DI3(mem_data_a_in[3]), 
        .DI4(mem_data_a_in[4]), .DI5(mem_data_a_in[5]), .DI6(mem_data_a_in[6]), 
        .DI7(mem_data_a_in[7]), .OE(net76341), .WEB(mem_we_a), .DO0(
        mem_data_a_out[0]), .DO1(mem_data_a_out[1]), .DO2(mem_data_a_out[2]), 
        .DO3(mem_data_a_out[3]), .DO4(mem_data_a_out[4]), .DO5(
        mem_data_a_out[5]), .DO6(mem_data_a_out[6]), .DO7(mem_data_a_out[7])
         );
  QDFFRBS mem_cs_a_reg ( .D(net76341), .CK(clk), .RB(n15893), .Q(mem_cs_a) );
  QDFFS image_size_in_reg_reg_1_ ( .D(image_size[1]), .CK(clk), .Q(
        image_size_in_reg[1]) );
  QDFFS image_size_in_reg_reg_0_ ( .D(image_size[0]), .CK(clk), .Q(
        image_size_in_reg[0]) );
  QDFFS action_in_reg_reg_2_ ( .D(action[2]), .CK(clk), .Q(action_in_reg[2])
         );
  QDFFS action_in_reg_reg_1_ ( .D(action[1]), .CK(clk), .Q(action_in_reg[1])
         );
  QDFFS action_in_reg_reg_0_ ( .D(action[0]), .CK(clk), .Q(action_in_reg[0])
         );
  QDFFS image_size_reg_master_reg_1_ ( .D(n15791), .CK(clk), .Q(
        image_size_reg_master[1]) );
  QDFFS image_size_reg_master_reg_0_ ( .D(n15790), .CK(clk), .Q(
        image_size_reg_master[0]) );
  QDFFS image_size_reg_set_reg_0_ ( .D(n15756), .CK(clk), .Q(
        image_size_reg_set[0]) );
  QDFFS medfilt_state_d1_reg_0_ ( .D(medfilt_state[0]), .CK(clk), .Q(
        medfilt_state_d1[0]) );
  QDFFS medfilt_cnt2_reg_0_ ( .D(n15736), .CK(clk), .Q(medfilt_cnt2[0]) );
  QDFFS medfilt_cnt2_d1_reg_0_ ( .D(medfilt_cnt2[0]), .CK(clk), .Q(
        medfilt_cnt2_d1[0]) );
  QDFFS medfilt_cnt2_reg_1_ ( .D(n15735), .CK(clk), .Q(medfilt_cnt2[1]) );
  QDFFS medfilt_cnt2_d1_reg_1_ ( .D(medfilt_cnt2[1]), .CK(clk), .Q(
        medfilt_cnt2_d1[1]) );
  QDFFS medfilt_cnt2_reg_2_ ( .D(n15734), .CK(clk), .Q(medfilt_cnt2[2]) );
  QDFFS medfilt_cnt2_d1_reg_2_ ( .D(medfilt_cnt2[2]), .CK(clk), .Q(
        medfilt_cnt2_d1[2]) );
  QDFFS medfilt_cnt2_reg_3_ ( .D(n15733), .CK(clk), .Q(medfilt_cnt2[3]) );
  QDFFS medfilt_cnt2_d1_reg_3_ ( .D(medfilt_cnt2[3]), .CK(clk), .Q(
        medfilt_cnt2_d1[3]) );
  QDFFS medfilt_state_d1_reg_2_ ( .D(medfilt_state[2]), .CK(clk), .Q(
        medfilt_state_d1[2]) );
  QDFFS action_done_reg ( .D(n15795), .CK(clk), .Q(action_done) );
  QDFFS action_reg_reg_7__0_ ( .D(n15788), .CK(clk), .Q(action_reg[21]) );
  QDFFS action_reg_reg_7__1_ ( .D(n15780), .CK(clk), .Q(action_reg[22]) );
  QDFFS action_reg_reg_7__2_ ( .D(n15772), .CK(clk), .Q(action_reg[23]) );
  QDFFS action_reg_reg_6__0_ ( .D(n15787), .CK(clk), .Q(action_reg[18]) );
  QDFFS action_reg_reg_5__0_ ( .D(n15786), .CK(clk), .Q(action_reg[15]) );
  QDFFS action_reg_reg_4__0_ ( .D(n15785), .CK(clk), .Q(action_reg[12]) );
  QDFFS action_reg_reg_3__0_ ( .D(n15784), .CK(clk), .Q(action_reg[9]) );
  QDFFS action_reg_reg_2__0_ ( .D(n15783), .CK(clk), .Q(action_reg[6]) );
  QDFFS action_reg_reg_1__0_ ( .D(n15782), .CK(clk), .Q(action_reg[3]) );
  QDFFS action_reg_reg_0__0_ ( .D(n15781), .CK(clk), .Q(action_reg[0]) );
  QDFFS action_reg_reg_6__1_ ( .D(n15779), .CK(clk), .Q(action_reg[19]) );
  QDFFS action_reg_reg_5__1_ ( .D(n15778), .CK(clk), .Q(action_reg[16]) );
  QDFFS action_reg_reg_4__1_ ( .D(n15777), .CK(clk), .Q(action_reg[13]) );
  QDFFS action_reg_reg_3__1_ ( .D(n15776), .CK(clk), .Q(action_reg[10]) );
  QDFFS action_reg_reg_2__1_ ( .D(n15775), .CK(clk), .Q(action_reg[7]) );
  QDFFS action_reg_reg_1__1_ ( .D(n15774), .CK(clk), .Q(action_reg[4]) );
  QDFFS action_reg_reg_0__1_ ( .D(n15773), .CK(clk), .Q(action_reg[1]) );
  QDFFS action_reg_reg_6__2_ ( .D(n15771), .CK(clk), .Q(action_reg[20]) );
  QDFFS action_reg_reg_5__2_ ( .D(n15770), .CK(clk), .Q(action_reg[17]) );
  QDFFS action_reg_reg_4__2_ ( .D(n15769), .CK(clk), .Q(action_reg[14]) );
  QDFFS action_reg_reg_3__2_ ( .D(n15768), .CK(clk), .Q(action_reg[11]) );
  QDFFS action_reg_reg_2__2_ ( .D(n15767), .CK(clk), .Q(action_reg[8]) );
  QDFFS action_reg_reg_1__2_ ( .D(n15766), .CK(clk), .Q(action_reg[5]) );
  QDFFS action_reg_reg_0__2_ ( .D(n15765), .CK(clk), .Q(action_reg[2]) );
  QDFFS image_size_reg_set_reg_1_ ( .D(n15757), .CK(clk), .Q(
        image_size_reg_set[1]) );
  QDFFS cnt_dyn_d1_reg_0_ ( .D(cnt_dyn[0]), .CK(clk), .Q(cnt_dyn_d1[0]) );
  QDFFS cnt_dyn_d1_reg_1_ ( .D(cnt_dyn[1]), .CK(clk), .Q(cnt_dyn_d1[1]) );
  QDFFS cnt_dyn_d1_reg_2_ ( .D(cnt_dyn[2]), .CK(clk), .Q(cnt_dyn_d1[2]) );
  QDFFS cnt_dyn_d1_reg_3_ ( .D(cnt_dyn[3]), .CK(clk), .Q(cnt_dyn_d1[3]) );
  QDFFS cnt_bdyn_d1_reg_3_ ( .D(cnt_bdyn[3]), .CK(clk), .Q(cnt_bdyn_d1[3]) );
  QDFFS cnt_bdyn_d1_reg_2_ ( .D(cnt_bdyn[2]), .CK(clk), .Q(cnt_bdyn_d1[2]) );
  QDFFS cnt_bdyn_d1_reg_1_ ( .D(cnt_bdyn[1]), .CK(clk), .Q(cnt_bdyn_d1[1]) );
  QDFFS cnt_bdyn_d1_reg_0_ ( .D(cnt_bdyn[0]), .CK(clk), .Q(cnt_bdyn_d1[0]) );
  QDFFS medfilt_state_d1_reg_3_ ( .D(medfilt_state[3]), .CK(clk), .Q(
        medfilt_state_d1[3]) );
  QDFFS medfilt_cnt_reg_0_ ( .D(N7502), .CK(clk), .Q(medfilt_cnt[0]) );
  QDFFS medfilt_cnt_d1_reg_0_ ( .D(medfilt_cnt[0]), .CK(clk), .Q(
        medfilt_cnt_d1[0]) );
  QDFFS medfilt_cnt_reg_1_ ( .D(N7503), .CK(clk), .Q(medfilt_cnt[1]) );
  QDFFS medfilt_cnt_d1_reg_1_ ( .D(medfilt_cnt[1]), .CK(clk), .Q(
        medfilt_cnt_d1[1]) );
  QDFFS medfilt_cnt_reg_2_ ( .D(N7504), .CK(clk), .Q(medfilt_cnt[2]) );
  QDFFS medfilt_cnt_d1_reg_2_ ( .D(medfilt_cnt[2]), .CK(clk), .Q(
        medfilt_cnt_d1[2]) );
  QDFFS medfilt_cnt_reg_3_ ( .D(N7505), .CK(clk), .Q(medfilt_cnt[3]) );
  QDFFS medfilt_cnt_d1_reg_3_ ( .D(medfilt_cnt[3]), .CK(clk), .Q(
        medfilt_cnt_d1[3]) );
  QDFFS medfilt_state_d1_reg_1_ ( .D(n30453), .CK(clk), .Q(medfilt_state_d1[1]) );
  QDFFS template_reg_reg_1__0__0_ ( .D(n15708), .CK(clk), .Q(template_reg[24])
         );
  QDFFS template_reg_reg_1__0__1_ ( .D(n15707), .CK(clk), .Q(template_reg[25])
         );
  QDFFS template_reg_reg_1__0__2_ ( .D(n15706), .CK(clk), .Q(template_reg[26])
         );
  QDFFS template_reg_reg_1__0__3_ ( .D(n15705), .CK(clk), .Q(template_reg[27])
         );
  QDFFS template_reg_reg_1__0__4_ ( .D(n15704), .CK(clk), .Q(template_reg[28])
         );
  QDFFS template_reg_reg_1__0__5_ ( .D(n15703), .CK(clk), .Q(template_reg[29])
         );
  QDFFS template_reg_reg_1__0__6_ ( .D(n15702), .CK(clk), .Q(template_reg[30])
         );
  QDFFS template_reg_reg_1__0__7_ ( .D(n15701), .CK(clk), .Q(template_reg[31])
         );
  QDFFS template_reg_reg_1__1__0_ ( .D(n15700), .CK(clk), .Q(template_reg[32])
         );
  QDFFS template_reg_reg_1__1__1_ ( .D(n15699), .CK(clk), .Q(template_reg[33])
         );
  QDFFS template_reg_reg_1__1__2_ ( .D(n15698), .CK(clk), .Q(template_reg[34])
         );
  QDFFS template_reg_reg_1__1__3_ ( .D(n15697), .CK(clk), .Q(template_reg[35])
         );
  QDFFS template_reg_reg_1__1__4_ ( .D(n15696), .CK(clk), .Q(template_reg[36])
         );
  QDFFS template_reg_reg_1__1__5_ ( .D(n15695), .CK(clk), .Q(template_reg[37])
         );
  QDFFS template_reg_reg_1__1__6_ ( .D(n15694), .CK(clk), .Q(template_reg[38])
         );
  QDFFS template_reg_reg_1__1__7_ ( .D(n15693), .CK(clk), .Q(template_reg[39])
         );
  QDFFS template_reg_reg_1__2__0_ ( .D(n15692), .CK(clk), .Q(template_reg[40])
         );
  QDFFS template_reg_reg_1__2__1_ ( .D(n15691), .CK(clk), .Q(template_reg[41])
         );
  QDFFS template_reg_reg_1__2__2_ ( .D(n15690), .CK(clk), .Q(template_reg[42])
         );
  QDFFS template_reg_reg_1__2__3_ ( .D(n15689), .CK(clk), .Q(template_reg[43])
         );
  QDFFS template_reg_reg_1__2__4_ ( .D(n15688), .CK(clk), .Q(template_reg[44])
         );
  QDFFS template_reg_reg_1__2__5_ ( .D(n15687), .CK(clk), .Q(template_reg[45])
         );
  QDFFS template_reg_reg_1__2__6_ ( .D(n15686), .CK(clk), .Q(template_reg[46])
         );
  QDFFS template_reg_reg_1__2__7_ ( .D(n15685), .CK(clk), .Q(template_reg[47])
         );
  QDFFS action_5_flag_reg ( .D(n13612), .CK(clk), .Q(action_5_flag) );
  QDFFS gray_img_reg_0__0__6_ ( .D(n15465), .CK(clk), .Q(gray_img[6]) );
  QDFFS mem_data_out_reg_shift_0_reg_0__6_ ( .D(n15809), .CK(clk), .Q(
        mem_data_out_reg_shift_0[6]) );
  QDFFS mem_data_out_reg_shift_0_reg_1__6_ ( .D(mem_data_out_reg_shift_0[6]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[14]) );
  QDFFS mem_data_out_reg_shift_0_reg_2__6_ ( .D(mem_data_out_reg_shift_0[14]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[22]) );
  QDFFS mem_data_out_reg_shift_0_reg_3__6_ ( .D(mem_data_out_reg_shift_0[22]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[30]) );
  QDFFS mem_data_out_reg_shift_0_reg_4__6_ ( .D(mem_data_out_reg_shift_0[30]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[38]) );
  QDFFS mem_data_out_reg_shift_0_reg_5__6_ ( .D(mem_data_out_reg_shift_0[38]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[46]) );
  QDFFS mem_data_out_reg_shift_0_reg_6__6_ ( .D(mem_data_out_reg_shift_0[46]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[54]) );
  QDFFS mem_data_out_reg_shift_0_reg_7__6_ ( .D(mem_data_out_reg_shift_0[54]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[62]) );
  QDFFS mem_data_out_reg_shift_0_reg_8__6_ ( .D(mem_data_out_reg_shift_0[62]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[70]) );
  QDFFS mem_data_out_reg_shift_0_reg_9__6_ ( .D(mem_data_out_reg_shift_0[70]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[78]) );
  QDFFS mem_data_out_reg_shift_0_reg_10__6_ ( .D(mem_data_out_reg_shift_0[78]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[86]) );
  QDFFS mem_data_out_reg_shift_0_reg_11__6_ ( .D(mem_data_out_reg_shift_0[86]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[94]) );
  QDFFS mem_data_out_reg_shift_0_reg_12__6_ ( .D(mem_data_out_reg_shift_0[94]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[102]) );
  QDFFS mem_data_out_reg_shift_0_reg_13__6_ ( .D(mem_data_out_reg_shift_0[102]), .CK(clk), .Q(mem_data_out_reg_shift_0[110]) );
  QDFFS mem_data_out_reg_shift_0_reg_14__6_ ( .D(mem_data_out_reg_shift_0[110]), .CK(clk), .Q(mem_data_out_reg_shift_0[118]) );
  QDFFS mem_data_out_reg_shift_0_reg_15__6_ ( .D(mem_data_out_reg_shift_0[118]), .CK(clk), .Q(mem_data_out_reg_shift_0[126]) );
  QDFFS mem_data_out_reg_shift_1_reg_0__6_ ( .D(n15826), .CK(clk), .Q(
        mem_data_out_reg_shift_1[6]) );
  QDFFS mem_data_out_reg_shift_1_reg_1__6_ ( .D(mem_data_out_reg_shift_1[6]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[14]) );
  QDFFS mem_data_out_reg_shift_1_reg_3__6_ ( .D(mem_data_out_reg_shift_1[22]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[30]) );
  QDFFS mem_data_out_reg_shift_1_reg_4__6_ ( .D(mem_data_out_reg_shift_1[30]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[38]) );
  QDFFS mem_data_out_reg_shift_1_reg_5__6_ ( .D(mem_data_out_reg_shift_1[38]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[46]) );
  QDFFS mem_data_out_reg_shift_1_reg_6__6_ ( .D(mem_data_out_reg_shift_1[46]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[54]) );
  QDFFS mem_data_out_reg_shift_1_reg_7__6_ ( .D(mem_data_out_reg_shift_1[54]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[62]) );
  QDFFS mem_data_out_reg_shift_1_reg_8__6_ ( .D(mem_data_out_reg_shift_1[62]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[70]) );
  QDFFS mem_data_out_reg_shift_1_reg_9__6_ ( .D(mem_data_out_reg_shift_1[70]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[78]) );
  QDFFS mem_data_out_reg_shift_1_reg_10__6_ ( .D(mem_data_out_reg_shift_1[78]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[86]) );
  QDFFS mem_data_out_reg_shift_1_reg_11__6_ ( .D(mem_data_out_reg_shift_1[86]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[94]) );
  QDFFS mem_data_out_reg_shift_1_reg_12__6_ ( .D(mem_data_out_reg_shift_1[94]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[102]) );
  QDFFS mem_data_out_reg_shift_1_reg_13__6_ ( .D(mem_data_out_reg_shift_1[102]), .CK(clk), .Q(mem_data_out_reg_shift_1[110]) );
  QDFFS mem_data_out_reg_shift_1_reg_14__6_ ( .D(mem_data_out_reg_shift_1[110]), .CK(clk), .Q(mem_data_out_reg_shift_1[118]) );
  QDFFS mem_data_out_reg_shift_1_reg_15__6_ ( .D(mem_data_out_reg_shift_1[118]), .CK(clk), .Q(mem_data_out_reg_shift_1[126]) );
  QDFFS mem_data_out_reg_shift_2_reg_0__6_ ( .D(n15834), .CK(clk), .Q(
        mem_data_out_reg_shift_2[6]) );
  QDFFS mem_data_out_reg_shift_2_reg_1__6_ ( .D(mem_data_out_reg_shift_2[6]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[14]) );
  QDFFS mem_data_out_reg_shift_2_reg_2__6_ ( .D(mem_data_out_reg_shift_2[14]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[22]) );
  QDFFS mem_data_out_reg_shift_2_reg_3__6_ ( .D(mem_data_out_reg_shift_2[22]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[30]) );
  QDFFS gray_img_reg_0__8__6_ ( .D(n15464), .CK(clk), .Q(gray_img[70]) );
  QDFFS gray_img_reg_0__9__6_ ( .D(n15463), .CK(clk), .Q(gray_img[78]) );
  QDFFS gray_img_reg_0__10__6_ ( .D(n15462), .CK(clk), .Q(gray_img[86]) );
  QDFFS gray_img_reg_0__11__6_ ( .D(n15461), .CK(clk), .Q(gray_img[94]) );
  QDFFS gray_img_reg_0__12__6_ ( .D(n15460), .CK(clk), .Q(gray_img[102]) );
  QDFFS gray_img_reg_0__13__6_ ( .D(n15459), .CK(clk), .Q(gray_img[110]) );
  QDFFS gray_img_reg_0__14__6_ ( .D(n15458), .CK(clk), .Q(gray_img[118]) );
  QDFFS gray_img_reg_0__15__6_ ( .D(n15457), .CK(clk), .Q(gray_img[126]) );
  QDFFS gray_img_reg_1__8__6_ ( .D(n15456), .CK(clk), .Q(gray_img[198]) );
  QDFFS gray_img_reg_1__9__6_ ( .D(n15455), .CK(clk), .Q(gray_img[206]) );
  QDFFS gray_img_reg_1__10__6_ ( .D(n15454), .CK(clk), .Q(gray_img[214]) );
  QDFFS gray_img_reg_1__11__6_ ( .D(n15453), .CK(clk), .Q(gray_img[222]) );
  QDFFS gray_img_reg_1__12__6_ ( .D(n15452), .CK(clk), .Q(gray_img[230]) );
  QDFFS gray_img_reg_1__13__6_ ( .D(n15451), .CK(clk), .Q(gray_img[238]) );
  QDFFS gray_img_reg_1__14__6_ ( .D(n15450), .CK(clk), .Q(gray_img[246]) );
  QDFFS gray_img_reg_1__15__6_ ( .D(n15449), .CK(clk), .Q(gray_img[254]) );
  QDFFS gray_img_reg_2__8__6_ ( .D(n15448), .CK(clk), .Q(gray_img[326]) );
  QDFFS gray_img_reg_2__9__6_ ( .D(n15447), .CK(clk), .Q(gray_img[334]) );
  QDFFS gray_img_reg_2__10__6_ ( .D(n15446), .CK(clk), .Q(gray_img[342]) );
  QDFFS gray_img_reg_2__11__6_ ( .D(n15445), .CK(clk), .Q(gray_img[350]) );
  QDFFS gray_img_reg_2__12__6_ ( .D(n15444), .CK(clk), .Q(gray_img[358]) );
  QDFFS gray_img_reg_2__13__6_ ( .D(n15443), .CK(clk), .Q(gray_img[366]) );
  QDFFS gray_img_reg_2__14__6_ ( .D(n15442), .CK(clk), .Q(gray_img[374]) );
  QDFFS gray_img_reg_2__15__6_ ( .D(n15441), .CK(clk), .Q(gray_img[382]) );
  QDFFS gray_img_reg_3__8__6_ ( .D(n15440), .CK(clk), .Q(gray_img[454]) );
  QDFFS gray_img_reg_3__9__6_ ( .D(n15439), .CK(clk), .Q(gray_img[462]) );
  QDFFS gray_img_reg_3__10__6_ ( .D(n15438), .CK(clk), .Q(gray_img[470]) );
  QDFFS gray_img_reg_3__11__6_ ( .D(n15437), .CK(clk), .Q(gray_img[478]) );
  QDFFS gray_img_reg_3__12__6_ ( .D(n15436), .CK(clk), .Q(gray_img[486]) );
  QDFFS gray_img_reg_3__13__6_ ( .D(n15435), .CK(clk), .Q(gray_img[494]) );
  QDFFS gray_img_reg_3__14__6_ ( .D(n15434), .CK(clk), .Q(gray_img[502]) );
  QDFFS gray_img_reg_3__15__6_ ( .D(n15433), .CK(clk), .Q(gray_img[510]) );
  QDFFS gray_img_reg_4__8__6_ ( .D(n15432), .CK(clk), .Q(gray_img[582]) );
  QDFFS gray_img_reg_4__9__6_ ( .D(n15431), .CK(clk), .Q(gray_img[590]) );
  QDFFS gray_img_reg_4__10__6_ ( .D(n15430), .CK(clk), .Q(gray_img[598]) );
  QDFFS gray_img_reg_4__11__6_ ( .D(n15429), .CK(clk), .Q(gray_img[606]) );
  QDFFS gray_img_reg_4__12__6_ ( .D(n15428), .CK(clk), .Q(gray_img[614]) );
  QDFFS gray_img_reg_4__13__6_ ( .D(n15427), .CK(clk), .Q(gray_img[622]) );
  QDFFS gray_img_reg_4__14__6_ ( .D(n15426), .CK(clk), .Q(gray_img[630]) );
  QDFFS gray_img_reg_4__15__6_ ( .D(n15425), .CK(clk), .Q(gray_img[638]) );
  QDFFS gray_img_reg_5__8__6_ ( .D(n15424), .CK(clk), .Q(gray_img[710]) );
  QDFFS gray_img_reg_5__9__6_ ( .D(n15423), .CK(clk), .Q(gray_img[718]) );
  QDFFS gray_img_reg_5__10__6_ ( .D(n15422), .CK(clk), .Q(gray_img[726]) );
  QDFFS gray_img_reg_5__11__6_ ( .D(n15421), .CK(clk), .Q(gray_img[734]) );
  QDFFS gray_img_reg_5__12__6_ ( .D(n15420), .CK(clk), .Q(gray_img[742]) );
  QDFFS gray_img_reg_5__13__6_ ( .D(n15419), .CK(clk), .Q(gray_img[750]) );
  QDFFS gray_img_reg_5__14__6_ ( .D(n15418), .CK(clk), .Q(gray_img[758]) );
  QDFFS gray_img_reg_5__15__6_ ( .D(n15417), .CK(clk), .Q(gray_img[766]) );
  QDFFS gray_img_reg_6__8__6_ ( .D(n15416), .CK(clk), .Q(gray_img[838]) );
  QDFFS gray_img_reg_6__9__6_ ( .D(n15415), .CK(clk), .Q(gray_img[846]) );
  QDFFS gray_img_reg_6__10__6_ ( .D(n15414), .CK(clk), .Q(gray_img[854]) );
  QDFFS gray_img_reg_6__11__6_ ( .D(n15413), .CK(clk), .Q(gray_img[862]) );
  QDFFS gray_img_reg_6__12__6_ ( .D(n15412), .CK(clk), .Q(gray_img[870]) );
  QDFFS gray_img_reg_6__13__6_ ( .D(n15411), .CK(clk), .Q(gray_img[878]) );
  QDFFS gray_img_reg_6__14__6_ ( .D(n15410), .CK(clk), .Q(gray_img[886]) );
  QDFFS gray_img_reg_6__15__6_ ( .D(n15409), .CK(clk), .Q(gray_img[894]) );
  QDFFS gray_img_reg_7__8__6_ ( .D(n15408), .CK(clk), .Q(gray_img[966]) );
  QDFFS gray_img_reg_7__9__6_ ( .D(n15407), .CK(clk), .Q(gray_img[974]) );
  QDFFS gray_img_reg_7__10__6_ ( .D(n15406), .CK(clk), .Q(gray_img[982]) );
  QDFFS gray_img_reg_7__11__6_ ( .D(n15405), .CK(clk), .Q(gray_img[990]) );
  QDFFS gray_img_reg_7__12__6_ ( .D(n15404), .CK(clk), .Q(gray_img[998]) );
  QDFFS gray_img_reg_7__13__6_ ( .D(n15403), .CK(clk), .Q(gray_img[1006]) );
  QDFFS gray_img_reg_7__14__6_ ( .D(n15402), .CK(clk), .Q(gray_img[1014]) );
  QDFFS gray_img_reg_7__15__6_ ( .D(n15401), .CK(clk), .Q(gray_img[1022]) );
  QDFFS gray_img_reg_8__0__6_ ( .D(n15400), .CK(clk), .Q(gray_img[1030]) );
  QDFFS gray_img_reg_8__1__6_ ( .D(n15399), .CK(clk), .Q(gray_img[1038]) );
  QDFFS gray_img_reg_8__2__6_ ( .D(n15398), .CK(clk), .Q(gray_img[1046]) );
  QDFFS gray_img_reg_8__3__6_ ( .D(n15397), .CK(clk), .Q(gray_img[1054]) );
  QDFFS gray_img_reg_8__4__6_ ( .D(n15396), .CK(clk), .Q(gray_img[1062]) );
  QDFFS gray_img_reg_8__5__6_ ( .D(n15395), .CK(clk), .Q(gray_img[1070]) );
  QDFFS gray_img_reg_8__6__6_ ( .D(n15394), .CK(clk), .Q(gray_img[1078]) );
  QDFFS gray_img_reg_8__7__6_ ( .D(n15393), .CK(clk), .Q(gray_img[1086]) );
  QDFFS gray_img_reg_8__8__6_ ( .D(n15392), .CK(clk), .Q(gray_img[1094]) );
  QDFFS gray_img_reg_8__9__6_ ( .D(n15391), .CK(clk), .Q(gray_img[1102]) );
  QDFFS gray_img_reg_8__10__6_ ( .D(n15390), .CK(clk), .Q(gray_img[1110]) );
  QDFFS gray_img_reg_8__11__6_ ( .D(n15389), .CK(clk), .Q(gray_img[1118]) );
  QDFFS gray_img_reg_8__12__6_ ( .D(n15388), .CK(clk), .Q(gray_img[1126]) );
  QDFFS gray_img_reg_8__13__6_ ( .D(n15387), .CK(clk), .Q(gray_img[1134]) );
  QDFFS gray_img_reg_8__14__6_ ( .D(n15386), .CK(clk), .Q(gray_img[1142]) );
  QDFFS gray_img_reg_8__15__6_ ( .D(n15385), .CK(clk), .Q(gray_img[1150]) );
  QDFFS gray_img_reg_9__0__6_ ( .D(n15384), .CK(clk), .Q(gray_img[1158]) );
  QDFFS gray_img_reg_9__1__6_ ( .D(n15383), .CK(clk), .Q(gray_img[1166]) );
  QDFFS gray_img_reg_9__2__6_ ( .D(n15382), .CK(clk), .Q(gray_img[1174]) );
  QDFFS gray_img_reg_9__3__6_ ( .D(n15381), .CK(clk), .Q(gray_img[1182]) );
  QDFFS gray_img_reg_9__4__6_ ( .D(n15380), .CK(clk), .Q(gray_img[1190]) );
  QDFFS gray_img_reg_9__5__6_ ( .D(n15379), .CK(clk), .Q(gray_img[1198]) );
  QDFFS gray_img_reg_9__6__6_ ( .D(n15378), .CK(clk), .Q(gray_img[1206]) );
  QDFFS gray_img_reg_9__7__6_ ( .D(n15377), .CK(clk), .Q(gray_img[1214]) );
  QDFFS gray_img_reg_9__8__6_ ( .D(n15376), .CK(clk), .Q(gray_img[1222]) );
  QDFFS gray_img_reg_9__9__6_ ( .D(n15375), .CK(clk), .Q(gray_img[1230]) );
  QDFFS gray_img_reg_9__10__6_ ( .D(n15374), .CK(clk), .Q(gray_img[1238]) );
  QDFFS gray_img_reg_9__11__6_ ( .D(n15373), .CK(clk), .Q(gray_img[1246]) );
  QDFFS gray_img_reg_9__12__6_ ( .D(n15372), .CK(clk), .Q(gray_img[1254]) );
  QDFFS gray_img_reg_9__13__6_ ( .D(n15371), .CK(clk), .Q(gray_img[1262]) );
  QDFFS gray_img_reg_9__14__6_ ( .D(n15370), .CK(clk), .Q(gray_img[1270]) );
  QDFFS gray_img_reg_9__15__6_ ( .D(n15369), .CK(clk), .Q(gray_img[1278]) );
  QDFFS gray_img_reg_10__0__6_ ( .D(n15368), .CK(clk), .Q(gray_img[1286]) );
  QDFFS gray_img_reg_10__1__6_ ( .D(n15367), .CK(clk), .Q(gray_img[1294]) );
  QDFFS gray_img_reg_10__2__6_ ( .D(n15366), .CK(clk), .Q(gray_img[1302]) );
  QDFFS gray_img_reg_10__3__6_ ( .D(n15365), .CK(clk), .Q(gray_img[1310]) );
  QDFFS gray_img_reg_10__4__6_ ( .D(n15364), .CK(clk), .Q(gray_img[1318]) );
  QDFFS gray_img_reg_10__5__6_ ( .D(n15363), .CK(clk), .Q(gray_img[1326]) );
  QDFFS gray_img_reg_10__6__6_ ( .D(n15362), .CK(clk), .Q(gray_img[1334]) );
  QDFFS gray_img_reg_10__7__6_ ( .D(n15361), .CK(clk), .Q(gray_img[1342]) );
  QDFFS gray_img_reg_10__8__6_ ( .D(n15360), .CK(clk), .Q(gray_img[1350]) );
  QDFFS gray_img_reg_10__9__6_ ( .D(n15359), .CK(clk), .Q(gray_img[1358]) );
  QDFFS gray_img_reg_10__10__6_ ( .D(n15358), .CK(clk), .Q(gray_img[1366]) );
  QDFFS gray_img_reg_10__11__6_ ( .D(n15357), .CK(clk), .Q(gray_img[1374]) );
  QDFFS gray_img_reg_10__12__6_ ( .D(n15356), .CK(clk), .Q(gray_img[1382]) );
  QDFFS gray_img_reg_10__13__6_ ( .D(n15355), .CK(clk), .Q(gray_img[1390]) );
  QDFFS gray_img_reg_10__14__6_ ( .D(n15354), .CK(clk), .Q(gray_img[1398]) );
  QDFFS gray_img_reg_10__15__6_ ( .D(n15353), .CK(clk), .Q(gray_img[1406]) );
  QDFFS gray_img_reg_11__0__6_ ( .D(n15352), .CK(clk), .Q(gray_img[1414]) );
  QDFFS gray_img_reg_11__1__6_ ( .D(n15351), .CK(clk), .Q(gray_img[1422]) );
  QDFFS gray_img_reg_11__2__6_ ( .D(n15350), .CK(clk), .Q(gray_img[1430]) );
  QDFFS gray_img_reg_11__3__6_ ( .D(n15349), .CK(clk), .Q(gray_img[1438]) );
  QDFFS gray_img_reg_11__4__6_ ( .D(n15348), .CK(clk), .Q(gray_img[1446]) );
  QDFFS gray_img_reg_11__5__6_ ( .D(n15347), .CK(clk), .Q(gray_img[1454]) );
  QDFFS gray_img_reg_11__6__6_ ( .D(n15346), .CK(clk), .Q(gray_img[1462]) );
  QDFFS gray_img_reg_11__7__6_ ( .D(n15345), .CK(clk), .Q(gray_img[1470]) );
  QDFFS gray_img_reg_11__8__6_ ( .D(n15344), .CK(clk), .Q(gray_img[1478]) );
  QDFFS gray_img_reg_11__9__6_ ( .D(n15343), .CK(clk), .Q(gray_img[1486]) );
  QDFFS gray_img_reg_11__10__6_ ( .D(n15342), .CK(clk), .Q(gray_img[1494]) );
  QDFFS gray_img_reg_11__11__6_ ( .D(n15341), .CK(clk), .Q(gray_img[1502]) );
  QDFFS gray_img_reg_11__12__6_ ( .D(n15340), .CK(clk), .Q(gray_img[1510]) );
  QDFFS gray_img_reg_11__13__6_ ( .D(n15339), .CK(clk), .Q(gray_img[1518]) );
  QDFFS gray_img_reg_11__14__6_ ( .D(n15338), .CK(clk), .Q(gray_img[1526]) );
  QDFFS gray_img_reg_11__15__6_ ( .D(n15337), .CK(clk), .Q(gray_img[1534]) );
  QDFFS gray_img_reg_12__0__6_ ( .D(n15336), .CK(clk), .Q(gray_img[1542]) );
  QDFFS gray_img_reg_12__1__6_ ( .D(n15335), .CK(clk), .Q(gray_img[1550]) );
  QDFFS gray_img_reg_12__2__6_ ( .D(n15334), .CK(clk), .Q(gray_img[1558]) );
  QDFFS gray_img_reg_12__3__6_ ( .D(n15333), .CK(clk), .Q(gray_img[1566]) );
  QDFFS gray_img_reg_12__4__6_ ( .D(n15332), .CK(clk), .Q(gray_img[1574]) );
  QDFFS gray_img_reg_12__5__6_ ( .D(n15331), .CK(clk), .Q(gray_img[1582]) );
  QDFFS gray_img_reg_12__6__6_ ( .D(n15330), .CK(clk), .Q(gray_img[1590]) );
  QDFFS gray_img_reg_12__7__6_ ( .D(n15329), .CK(clk), .Q(gray_img[1598]) );
  QDFFS gray_img_reg_12__8__6_ ( .D(n15328), .CK(clk), .Q(gray_img[1606]) );
  QDFFS gray_img_reg_12__9__6_ ( .D(n15327), .CK(clk), .Q(gray_img[1614]) );
  QDFFS gray_img_reg_12__10__6_ ( .D(n15326), .CK(clk), .Q(gray_img[1622]) );
  QDFFS gray_img_reg_12__11__6_ ( .D(n15325), .CK(clk), .Q(gray_img[1630]) );
  QDFFS gray_img_reg_12__12__6_ ( .D(n15324), .CK(clk), .Q(gray_img[1638]) );
  QDFFS gray_img_reg_12__13__6_ ( .D(n15323), .CK(clk), .Q(gray_img[1646]) );
  QDFFS gray_img_reg_12__14__6_ ( .D(n15322), .CK(clk), .Q(gray_img[1654]) );
  QDFFS gray_img_reg_12__15__6_ ( .D(n15321), .CK(clk), .Q(gray_img[1662]) );
  QDFFS gray_img_reg_13__0__6_ ( .D(n15320), .CK(clk), .Q(gray_img[1670]) );
  QDFFS gray_img_reg_13__1__6_ ( .D(n15319), .CK(clk), .Q(gray_img[1678]) );
  QDFFS gray_img_reg_13__2__6_ ( .D(n15318), .CK(clk), .Q(gray_img[1686]) );
  QDFFS gray_img_reg_13__3__6_ ( .D(n15317), .CK(clk), .Q(gray_img[1694]) );
  QDFFS gray_img_reg_13__4__6_ ( .D(n15316), .CK(clk), .Q(gray_img[1702]) );
  QDFFS gray_img_reg_13__5__6_ ( .D(n15315), .CK(clk), .Q(gray_img[1710]) );
  QDFFS gray_img_reg_13__6__6_ ( .D(n15314), .CK(clk), .Q(gray_img[1718]) );
  QDFFS gray_img_reg_13__7__6_ ( .D(n15313), .CK(clk), .Q(gray_img[1726]) );
  QDFFS gray_img_reg_13__8__6_ ( .D(n15312), .CK(clk), .Q(gray_img[1734]) );
  QDFFS gray_img_reg_13__9__6_ ( .D(n15311), .CK(clk), .Q(gray_img[1742]) );
  QDFFS gray_img_reg_13__10__6_ ( .D(n15310), .CK(clk), .Q(gray_img[1750]) );
  QDFFS gray_img_reg_13__11__6_ ( .D(n15309), .CK(clk), .Q(gray_img[1758]) );
  QDFFS gray_img_reg_13__12__6_ ( .D(n15308), .CK(clk), .Q(gray_img[1766]) );
  QDFFS gray_img_reg_13__13__6_ ( .D(n15307), .CK(clk), .Q(gray_img[1774]) );
  QDFFS gray_img_reg_13__14__6_ ( .D(n15306), .CK(clk), .Q(gray_img[1782]) );
  QDFFS gray_img_reg_13__15__6_ ( .D(n15305), .CK(clk), .Q(gray_img[1790]) );
  QDFFS gray_img_reg_14__0__6_ ( .D(n15304), .CK(clk), .Q(gray_img[1798]) );
  QDFFS gray_img_reg_14__1__6_ ( .D(n15303), .CK(clk), .Q(gray_img[1806]) );
  QDFFS gray_img_reg_14__2__6_ ( .D(n15302), .CK(clk), .Q(gray_img[1814]) );
  QDFFS gray_img_reg_14__3__6_ ( .D(n15301), .CK(clk), .Q(gray_img[1822]) );
  QDFFS gray_img_reg_14__4__6_ ( .D(n15300), .CK(clk), .Q(gray_img[1830]) );
  QDFFS gray_img_reg_14__5__6_ ( .D(n15299), .CK(clk), .Q(gray_img[1838]) );
  QDFFS gray_img_reg_14__6__6_ ( .D(n15298), .CK(clk), .Q(gray_img[1846]) );
  QDFFS gray_img_reg_14__7__6_ ( .D(n15297), .CK(clk), .Q(gray_img[1854]) );
  QDFFS gray_img_reg_14__8__6_ ( .D(n15296), .CK(clk), .Q(gray_img[1862]) );
  QDFFS gray_img_reg_14__9__6_ ( .D(n15295), .CK(clk), .Q(gray_img[1870]) );
  QDFFS gray_img_reg_14__10__6_ ( .D(n15294), .CK(clk), .Q(gray_img[1878]) );
  QDFFS gray_img_reg_14__11__6_ ( .D(n15293), .CK(clk), .Q(gray_img[1886]) );
  QDFFS gray_img_reg_14__12__6_ ( .D(n15292), .CK(clk), .Q(gray_img[1894]) );
  QDFFS gray_img_reg_14__13__6_ ( .D(n15291), .CK(clk), .Q(gray_img[1902]) );
  QDFFS gray_img_reg_14__14__6_ ( .D(n15290), .CK(clk), .Q(gray_img[1910]) );
  QDFFS gray_img_reg_14__15__6_ ( .D(n15289), .CK(clk), .Q(gray_img[1918]) );
  QDFFS gray_img_reg_15__0__6_ ( .D(n15288), .CK(clk), .Q(gray_img[1926]) );
  QDFFS gray_img_reg_15__1__6_ ( .D(n15287), .CK(clk), .Q(gray_img[1934]) );
  QDFFS gray_img_reg_15__2__6_ ( .D(n15286), .CK(clk), .Q(gray_img[1942]) );
  QDFFS gray_img_reg_15__3__6_ ( .D(n15285), .CK(clk), .Q(gray_img[1950]) );
  QDFFS gray_img_reg_15__4__6_ ( .D(n15284), .CK(clk), .Q(gray_img[1958]) );
  QDFFS gray_img_reg_15__5__6_ ( .D(n15283), .CK(clk), .Q(gray_img[1966]) );
  QDFFS gray_img_reg_15__6__6_ ( .D(n15282), .CK(clk), .Q(gray_img[1974]) );
  QDFFS gray_img_reg_15__7__6_ ( .D(n15281), .CK(clk), .Q(gray_img[1982]) );
  QDFFS gray_img_reg_15__8__6_ ( .D(n15280), .CK(clk), .Q(gray_img[1990]) );
  QDFFS gray_img_reg_15__9__6_ ( .D(n15279), .CK(clk), .Q(gray_img[1998]) );
  QDFFS gray_img_reg_15__10__6_ ( .D(n15278), .CK(clk), .Q(gray_img[2006]) );
  QDFFS gray_img_reg_15__11__6_ ( .D(n15277), .CK(clk), .Q(gray_img[2014]) );
  QDFFS gray_img_reg_15__12__6_ ( .D(n15276), .CK(clk), .Q(gray_img[2022]) );
  QDFFS gray_img_reg_15__13__6_ ( .D(n15275), .CK(clk), .Q(gray_img[2030]) );
  QDFFS gray_img_reg_15__14__6_ ( .D(n15274), .CK(clk), .Q(gray_img[2038]) );
  QDFFS gray_img_reg_15__15__6_ ( .D(n15273), .CK(clk), .Q(gray_img[2046]) );
  QDFFS gray_img_reg_7__5__6_ ( .D(n15270), .CK(clk), .Q(gray_img[942]) );
  QDFFS gray_img_reg_0__4__6_ ( .D(n14251), .CK(clk), .Q(gray_img[38]) );
  QDFFS gray_img_reg_0__5__6_ ( .D(n14242), .CK(clk), .Q(gray_img[46]) );
  QDFFS gray_img_reg_0__6__6_ ( .D(n14233), .CK(clk), .Q(gray_img[54]) );
  QDFFS gray_img_reg_0__7__6_ ( .D(n14224), .CK(clk), .Q(gray_img[62]) );
  QDFFS gray_img_reg_1__4__6_ ( .D(n14207), .CK(clk), .Q(gray_img[166]) );
  QDFFS gray_img_reg_1__5__6_ ( .D(n14198), .CK(clk), .Q(gray_img[174]) );
  QDFFS gray_img_reg_1__6__6_ ( .D(n14189), .CK(clk), .Q(gray_img[182]) );
  QDFFS gray_img_reg_1__7__6_ ( .D(n14180), .CK(clk), .Q(gray_img[190]) );
  QDFFS gray_img_reg_2__4__6_ ( .D(n14163), .CK(clk), .Q(gray_img[294]) );
  QDFFS gray_img_reg_2__5__6_ ( .D(n14154), .CK(clk), .Q(gray_img[302]) );
  QDFFS gray_img_reg_2__6__6_ ( .D(n14145), .CK(clk), .Q(gray_img[310]) );
  QDFFS gray_img_reg_2__7__6_ ( .D(n14136), .CK(clk), .Q(gray_img[318]) );
  QDFFS gray_img_reg_3__4__6_ ( .D(n14119), .CK(clk), .Q(gray_img[422]) );
  QDFFS gray_img_reg_3__5__6_ ( .D(n14110), .CK(clk), .Q(gray_img[430]) );
  QDFFS gray_img_reg_3__6__6_ ( .D(n14101), .CK(clk), .Q(gray_img[438]) );
  QDFFS gray_img_reg_3__7__6_ ( .D(n14092), .CK(clk), .Q(gray_img[446]) );
  QDFFS gray_img_reg_4__0__6_ ( .D(n14067), .CK(clk), .Q(gray_img[518]) );
  QDFFS gray_img_reg_4__1__6_ ( .D(n14058), .CK(clk), .Q(gray_img[526]) );
  QDFFS gray_img_reg_4__2__6_ ( .D(n14049), .CK(clk), .Q(gray_img[534]) );
  QDFFS gray_img_reg_4__3__6_ ( .D(n14040), .CK(clk), .Q(gray_img[542]) );
  QDFFS gray_img_reg_4__4__6_ ( .D(n14031), .CK(clk), .Q(gray_img[550]) );
  QDFFS gray_img_reg_4__5__6_ ( .D(n14022), .CK(clk), .Q(gray_img[558]) );
  QDFFS gray_img_reg_4__6__6_ ( .D(n14013), .CK(clk), .Q(gray_img[566]) );
  QDFFS gray_img_reg_4__7__6_ ( .D(n14004), .CK(clk), .Q(gray_img[574]) );
  QDFFS gray_img_reg_5__0__6_ ( .D(n13979), .CK(clk), .Q(gray_img[646]) );
  QDFFS gray_img_reg_5__1__6_ ( .D(n13970), .CK(clk), .Q(gray_img[654]) );
  QDFFS gray_img_reg_5__2__6_ ( .D(n13961), .CK(clk), .Q(gray_img[662]) );
  QDFFS gray_img_reg_5__3__6_ ( .D(n13953), .CK(clk), .Q(gray_img[670]) );
  QDFFS gray_img_reg_5__4__6_ ( .D(n13945), .CK(clk), .Q(gray_img[678]) );
  QDFFS gray_img_reg_5__5__6_ ( .D(n13938), .CK(clk), .Q(gray_img[686]) );
  QDFFS gray_img_reg_5__6__6_ ( .D(n13931), .CK(clk), .Q(gray_img[694]) );
  QDFFS gray_img_reg_5__7__6_ ( .D(n13925), .CK(clk), .Q(gray_img[702]) );
  QDFFS gray_img_reg_6__0__6_ ( .D(n13903), .CK(clk), .Q(gray_img[774]) );
  QDFFS gray_img_reg_6__1__6_ ( .D(n13897), .CK(clk), .Q(gray_img[782]) );
  QDFFS gray_img_reg_6__2__6_ ( .D(n13891), .CK(clk), .Q(gray_img[790]) );
  QDFFS gray_img_reg_6__3__6_ ( .D(n13885), .CK(clk), .Q(gray_img[798]) );
  QDFFS gray_img_reg_6__4__6_ ( .D(n13879), .CK(clk), .Q(gray_img[806]) );
  QDFFS gray_img_reg_6__5__6_ ( .D(n13873), .CK(clk), .Q(gray_img[814]) );
  QDFFS gray_img_reg_6__6__6_ ( .D(n13867), .CK(clk), .Q(gray_img[822]) );
  QDFFS gray_img_reg_6__7__6_ ( .D(n13861), .CK(clk), .Q(gray_img[830]) );
  QDFFS gray_img_reg_7__0__6_ ( .D(n13839), .CK(clk), .Q(gray_img[902]) );
  QDFFS gray_img_reg_7__1__6_ ( .D(n13834), .CK(clk), .Q(gray_img[910]) );
  QDFFS gray_img_reg_7__2__6_ ( .D(n13829), .CK(clk), .Q(gray_img[918]) );
  QDFFS gray_img_reg_7__3__6_ ( .D(n13825), .CK(clk), .Q(gray_img[926]) );
  QDFFS gray_img_reg_3__1__6_ ( .D(n15071), .CK(clk), .Q(gray_img[398]) );
  QDFFS gray_img_reg_7__4__6_ ( .D(n13821), .CK(clk), .Q(gray_img[934]) );
  QDFFS gray_img_reg_0__2__6_ ( .D(n13796), .CK(clk), .Q(gray_img[22]) );
  QDFFS gray_img_reg_0__3__6_ ( .D(n13786), .CK(clk), .Q(gray_img[30]) );
  QDFFS gray_img_reg_1__2__6_ ( .D(n13766), .CK(clk), .Q(gray_img[150]) );
  QDFFS gray_img_reg_1__3__6_ ( .D(n13756), .CK(clk), .Q(gray_img[158]) );
  QDFFS gray_img_reg_0__1__6_ ( .D(n13748), .CK(clk), .Q(gray_img[14]) );
  QDFFS gray_img_reg_2__0__6_ ( .D(n13730), .CK(clk), .Q(gray_img[262]) );
  QDFFS gray_img_reg_2__1__6_ ( .D(n13701), .CK(clk), .Q(gray_img[270]) );
  QDFFS gray_img_reg_2__2__6_ ( .D(n13675), .CK(clk), .Q(gray_img[278]) );
  QDFFS gray_img_reg_2__3__6_ ( .D(n13652), .CK(clk), .Q(gray_img[286]) );
  QDFFS gray_img_reg_3__0__6_ ( .D(n13632), .CK(clk), .Q(gray_img[390]) );
  QDFFS gray_img_reg_1__0__6_ ( .D(n13623), .CK(clk), .Q(gray_img[134]) );
  QDFFS gray_img_reg_3__2__6_ ( .D(n13617), .CK(clk), .Q(gray_img[406]) );
  QDFFS gray_img_reg_7__6__6_ ( .D(n13615), .CK(clk), .Q(gray_img[950]) );
  QDFFS gray_img_reg_7__7__6_ ( .D(n13614), .CK(clk), .Q(gray_img[958]) );
  QDFFS gray_img_reg_3__3__6_ ( .D(n15271), .CK(clk), .Q(gray_img[414]) );
  QDFFS gray_img_reg_1__1__6_ ( .D(n15272), .CK(clk), .Q(gray_img[142]) );
  QDFFS gray_img_reg_0__0__5_ ( .D(n15076), .CK(clk), .Q(gray_img[5]) );
  QDFFS mem_data_out_reg_shift_0_reg_0__5_ ( .D(n15810), .CK(clk), .Q(
        mem_data_out_reg_shift_0[5]) );
  QDFFS mem_data_out_reg_shift_0_reg_1__5_ ( .D(mem_data_out_reg_shift_0[5]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[13]) );
  QDFFS mem_data_out_reg_shift_0_reg_2__5_ ( .D(mem_data_out_reg_shift_0[13]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[21]) );
  QDFFS mem_data_out_reg_shift_0_reg_3__5_ ( .D(mem_data_out_reg_shift_0[21]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[29]) );
  QDFFS mem_data_out_reg_shift_0_reg_4__5_ ( .D(mem_data_out_reg_shift_0[29]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[37]) );
  QDFFS mem_data_out_reg_shift_0_reg_5__5_ ( .D(mem_data_out_reg_shift_0[37]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[45]) );
  QDFFS mem_data_out_reg_shift_0_reg_6__5_ ( .D(mem_data_out_reg_shift_0[45]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[53]) );
  QDFFS mem_data_out_reg_shift_0_reg_7__5_ ( .D(mem_data_out_reg_shift_0[53]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[61]) );
  QDFFS mem_data_out_reg_shift_0_reg_8__5_ ( .D(mem_data_out_reg_shift_0[61]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[69]) );
  QDFFS mem_data_out_reg_shift_0_reg_9__5_ ( .D(mem_data_out_reg_shift_0[69]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[77]) );
  QDFFS mem_data_out_reg_shift_0_reg_10__5_ ( .D(mem_data_out_reg_shift_0[77]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[85]) );
  QDFFS mem_data_out_reg_shift_0_reg_11__5_ ( .D(mem_data_out_reg_shift_0[85]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[93]) );
  QDFFS mem_data_out_reg_shift_0_reg_12__5_ ( .D(mem_data_out_reg_shift_0[93]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[101]) );
  QDFFS mem_data_out_reg_shift_0_reg_13__5_ ( .D(mem_data_out_reg_shift_0[101]), .CK(clk), .Q(mem_data_out_reg_shift_0[109]) );
  QDFFS mem_data_out_reg_shift_0_reg_14__5_ ( .D(mem_data_out_reg_shift_0[109]), .CK(clk), .Q(mem_data_out_reg_shift_0[117]) );
  QDFFS mem_data_out_reg_shift_0_reg_15__5_ ( .D(mem_data_out_reg_shift_0[117]), .CK(clk), .Q(mem_data_out_reg_shift_0[125]) );
  QDFFS mem_data_out_reg_shift_1_reg_0__5_ ( .D(n15827), .CK(clk), .Q(
        mem_data_out_reg_shift_1[5]) );
  QDFFS mem_data_out_reg_shift_1_reg_1__5_ ( .D(mem_data_out_reg_shift_1[5]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[13]) );
  QDFFS mem_data_out_reg_shift_1_reg_3__5_ ( .D(mem_data_out_reg_shift_1[21]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[29]) );
  QDFFS mem_data_out_reg_shift_1_reg_4__5_ ( .D(mem_data_out_reg_shift_1[29]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[37]) );
  QDFFS mem_data_out_reg_shift_1_reg_5__5_ ( .D(mem_data_out_reg_shift_1[37]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[45]) );
  QDFFS mem_data_out_reg_shift_1_reg_6__5_ ( .D(mem_data_out_reg_shift_1[45]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[53]) );
  QDFFS mem_data_out_reg_shift_1_reg_7__5_ ( .D(mem_data_out_reg_shift_1[53]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[61]) );
  QDFFS mem_data_out_reg_shift_1_reg_8__5_ ( .D(mem_data_out_reg_shift_1[61]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[69]) );
  QDFFS mem_data_out_reg_shift_1_reg_9__5_ ( .D(mem_data_out_reg_shift_1[69]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[77]) );
  QDFFS mem_data_out_reg_shift_1_reg_10__5_ ( .D(mem_data_out_reg_shift_1[77]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[85]) );
  QDFFS mem_data_out_reg_shift_1_reg_11__5_ ( .D(mem_data_out_reg_shift_1[85]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[93]) );
  QDFFS mem_data_out_reg_shift_1_reg_12__5_ ( .D(mem_data_out_reg_shift_1[93]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[101]) );
  QDFFS mem_data_out_reg_shift_1_reg_13__5_ ( .D(mem_data_out_reg_shift_1[101]), .CK(clk), .Q(mem_data_out_reg_shift_1[109]) );
  QDFFS mem_data_out_reg_shift_1_reg_14__5_ ( .D(mem_data_out_reg_shift_1[109]), .CK(clk), .Q(mem_data_out_reg_shift_1[117]) );
  QDFFS mem_data_out_reg_shift_1_reg_15__5_ ( .D(mem_data_out_reg_shift_1[117]), .CK(clk), .Q(mem_data_out_reg_shift_1[125]) );
  QDFFS mem_data_out_reg_shift_2_reg_0__5_ ( .D(n15835), .CK(clk), .Q(
        mem_data_out_reg_shift_2[5]) );
  QDFFS mem_data_out_reg_shift_2_reg_1__5_ ( .D(mem_data_out_reg_shift_2[5]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[13]) );
  QDFFS mem_data_out_reg_shift_2_reg_2__5_ ( .D(mem_data_out_reg_shift_2[13]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[21]) );
  QDFFS mem_data_out_reg_shift_2_reg_3__5_ ( .D(mem_data_out_reg_shift_2[21]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[29]) );
  QDFFS gray_img_reg_0__8__5_ ( .D(n15268), .CK(clk), .Q(gray_img[69]) );
  QDFFS gray_img_reg_0__9__5_ ( .D(n15267), .CK(clk), .Q(gray_img[77]) );
  QDFFS gray_img_reg_0__10__5_ ( .D(n15266), .CK(clk), .Q(gray_img[85]) );
  QDFFS gray_img_reg_0__11__5_ ( .D(n15265), .CK(clk), .Q(gray_img[93]) );
  QDFFS gray_img_reg_0__12__5_ ( .D(n15264), .CK(clk), .Q(gray_img[101]) );
  QDFFS gray_img_reg_0__13__5_ ( .D(n15263), .CK(clk), .Q(gray_img[109]) );
  QDFFS gray_img_reg_0__14__5_ ( .D(n15262), .CK(clk), .Q(gray_img[117]) );
  QDFFS gray_img_reg_0__15__5_ ( .D(n15261), .CK(clk), .Q(gray_img[125]) );
  QDFFS gray_img_reg_1__8__5_ ( .D(n15260), .CK(clk), .Q(gray_img[197]) );
  QDFFS gray_img_reg_1__9__5_ ( .D(n15259), .CK(clk), .Q(gray_img[205]) );
  QDFFS gray_img_reg_1__10__5_ ( .D(n15258), .CK(clk), .Q(gray_img[213]) );
  QDFFS gray_img_reg_1__11__5_ ( .D(n15257), .CK(clk), .Q(gray_img[221]) );
  QDFFS gray_img_reg_1__12__5_ ( .D(n15256), .CK(clk), .Q(gray_img[229]) );
  QDFFS gray_img_reg_1__13__5_ ( .D(n15255), .CK(clk), .Q(gray_img[237]) );
  QDFFS gray_img_reg_1__14__5_ ( .D(n15254), .CK(clk), .Q(gray_img[245]) );
  QDFFS gray_img_reg_1__15__5_ ( .D(n15253), .CK(clk), .Q(gray_img[253]) );
  QDFFS gray_img_reg_2__8__5_ ( .D(n15252), .CK(clk), .Q(gray_img[325]) );
  QDFFS gray_img_reg_2__9__5_ ( .D(n15251), .CK(clk), .Q(gray_img[333]) );
  QDFFS gray_img_reg_2__10__5_ ( .D(n15250), .CK(clk), .Q(gray_img[341]) );
  QDFFS gray_img_reg_2__11__5_ ( .D(n15249), .CK(clk), .Q(gray_img[349]) );
  QDFFS gray_img_reg_2__12__5_ ( .D(n15248), .CK(clk), .Q(gray_img[357]) );
  QDFFS gray_img_reg_2__13__5_ ( .D(n15247), .CK(clk), .Q(gray_img[365]) );
  QDFFS gray_img_reg_2__14__5_ ( .D(n15246), .CK(clk), .Q(gray_img[373]) );
  QDFFS gray_img_reg_2__15__5_ ( .D(n15245), .CK(clk), .Q(gray_img[381]) );
  QDFFS gray_img_reg_3__8__5_ ( .D(n15244), .CK(clk), .Q(gray_img[453]) );
  QDFFS gray_img_reg_3__9__5_ ( .D(n15243), .CK(clk), .Q(gray_img[461]) );
  QDFFS gray_img_reg_3__10__5_ ( .D(n15242), .CK(clk), .Q(gray_img[469]) );
  QDFFS gray_img_reg_3__11__5_ ( .D(n15241), .CK(clk), .Q(gray_img[477]) );
  QDFFS gray_img_reg_3__12__5_ ( .D(n15240), .CK(clk), .Q(gray_img[485]) );
  QDFFS gray_img_reg_3__13__5_ ( .D(n15239), .CK(clk), .Q(gray_img[493]) );
  QDFFS gray_img_reg_3__14__5_ ( .D(n15238), .CK(clk), .Q(gray_img[501]) );
  QDFFS gray_img_reg_3__15__5_ ( .D(n15237), .CK(clk), .Q(gray_img[509]) );
  QDFFS gray_img_reg_4__8__5_ ( .D(n15236), .CK(clk), .Q(gray_img[581]) );
  QDFFS gray_img_reg_4__9__5_ ( .D(n15235), .CK(clk), .Q(gray_img[589]) );
  QDFFS gray_img_reg_4__10__5_ ( .D(n15234), .CK(clk), .Q(gray_img[597]) );
  QDFFS gray_img_reg_4__11__5_ ( .D(n15233), .CK(clk), .Q(gray_img[605]) );
  QDFFS gray_img_reg_4__12__5_ ( .D(n15232), .CK(clk), .Q(gray_img[613]) );
  QDFFS gray_img_reg_4__13__5_ ( .D(n15231), .CK(clk), .Q(gray_img[621]) );
  QDFFS gray_img_reg_4__14__5_ ( .D(n15230), .CK(clk), .Q(gray_img[629]) );
  QDFFS gray_img_reg_4__15__5_ ( .D(n15229), .CK(clk), .Q(gray_img[637]) );
  QDFFS gray_img_reg_5__8__5_ ( .D(n15228), .CK(clk), .Q(gray_img[709]) );
  QDFFS gray_img_reg_5__9__5_ ( .D(n15227), .CK(clk), .Q(gray_img[717]) );
  QDFFS gray_img_reg_5__10__5_ ( .D(n15226), .CK(clk), .Q(gray_img[725]) );
  QDFFS gray_img_reg_5__11__5_ ( .D(n15225), .CK(clk), .Q(gray_img[733]) );
  QDFFS gray_img_reg_5__12__5_ ( .D(n15224), .CK(clk), .Q(gray_img[741]) );
  QDFFS gray_img_reg_5__13__5_ ( .D(n15223), .CK(clk), .Q(gray_img[749]) );
  QDFFS gray_img_reg_5__14__5_ ( .D(n15222), .CK(clk), .Q(gray_img[757]) );
  QDFFS gray_img_reg_5__15__5_ ( .D(n15221), .CK(clk), .Q(gray_img[765]) );
  QDFFS gray_img_reg_6__8__5_ ( .D(n15220), .CK(clk), .Q(gray_img[837]) );
  QDFFS gray_img_reg_6__9__5_ ( .D(n15219), .CK(clk), .Q(gray_img[845]) );
  QDFFS gray_img_reg_6__10__5_ ( .D(n15218), .CK(clk), .Q(gray_img[853]) );
  QDFFS gray_img_reg_6__11__5_ ( .D(n15217), .CK(clk), .Q(gray_img[861]) );
  QDFFS gray_img_reg_6__12__5_ ( .D(n15216), .CK(clk), .Q(gray_img[869]) );
  QDFFS gray_img_reg_6__13__5_ ( .D(n15215), .CK(clk), .Q(gray_img[877]) );
  QDFFS gray_img_reg_6__14__5_ ( .D(n15214), .CK(clk), .Q(gray_img[885]) );
  QDFFS gray_img_reg_6__15__5_ ( .D(n15213), .CK(clk), .Q(gray_img[893]) );
  QDFFS gray_img_reg_7__8__5_ ( .D(n15212), .CK(clk), .Q(gray_img[965]) );
  QDFFS gray_img_reg_7__9__5_ ( .D(n15211), .CK(clk), .Q(gray_img[973]) );
  QDFFS gray_img_reg_7__10__5_ ( .D(n15210), .CK(clk), .Q(gray_img[981]) );
  QDFFS gray_img_reg_7__11__5_ ( .D(n15209), .CK(clk), .Q(gray_img[989]) );
  QDFFS gray_img_reg_7__12__5_ ( .D(n15208), .CK(clk), .Q(gray_img[997]) );
  QDFFS gray_img_reg_7__13__5_ ( .D(n15207), .CK(clk), .Q(gray_img[1005]) );
  QDFFS gray_img_reg_7__14__5_ ( .D(n15206), .CK(clk), .Q(gray_img[1013]) );
  QDFFS gray_img_reg_7__15__5_ ( .D(n15205), .CK(clk), .Q(gray_img[1021]) );
  QDFFS gray_img_reg_8__0__5_ ( .D(n15204), .CK(clk), .Q(gray_img[1029]) );
  QDFFS gray_img_reg_8__1__5_ ( .D(n15203), .CK(clk), .Q(gray_img[1037]) );
  QDFFS gray_img_reg_8__2__5_ ( .D(n15202), .CK(clk), .Q(gray_img[1045]) );
  QDFFS gray_img_reg_8__3__5_ ( .D(n15201), .CK(clk), .Q(gray_img[1053]) );
  QDFFS gray_img_reg_8__4__5_ ( .D(n15200), .CK(clk), .Q(gray_img[1061]) );
  QDFFS gray_img_reg_8__5__5_ ( .D(n15199), .CK(clk), .Q(gray_img[1069]) );
  QDFFS gray_img_reg_8__6__5_ ( .D(n15198), .CK(clk), .Q(gray_img[1077]) );
  QDFFS gray_img_reg_8__7__5_ ( .D(n15197), .CK(clk), .Q(gray_img[1085]) );
  QDFFS gray_img_reg_8__8__5_ ( .D(n15196), .CK(clk), .Q(gray_img[1093]) );
  QDFFS gray_img_reg_8__9__5_ ( .D(n15195), .CK(clk), .Q(gray_img[1101]) );
  QDFFS gray_img_reg_8__10__5_ ( .D(n15194), .CK(clk), .Q(gray_img[1109]) );
  QDFFS gray_img_reg_8__11__5_ ( .D(n15193), .CK(clk), .Q(gray_img[1117]) );
  QDFFS gray_img_reg_8__12__5_ ( .D(n15192), .CK(clk), .Q(gray_img[1125]) );
  QDFFS gray_img_reg_8__13__5_ ( .D(n15191), .CK(clk), .Q(gray_img[1133]) );
  QDFFS gray_img_reg_8__14__5_ ( .D(n15190), .CK(clk), .Q(gray_img[1141]) );
  QDFFS gray_img_reg_8__15__5_ ( .D(n15189), .CK(clk), .Q(gray_img[1149]) );
  QDFFS gray_img_reg_9__0__5_ ( .D(n15188), .CK(clk), .Q(gray_img[1157]) );
  QDFFS gray_img_reg_9__1__5_ ( .D(n15187), .CK(clk), .Q(gray_img[1165]) );
  QDFFS gray_img_reg_9__2__5_ ( .D(n15186), .CK(clk), .Q(gray_img[1173]) );
  QDFFS gray_img_reg_9__3__5_ ( .D(n15185), .CK(clk), .Q(gray_img[1181]) );
  QDFFS gray_img_reg_9__4__5_ ( .D(n15184), .CK(clk), .Q(gray_img[1189]) );
  QDFFS gray_img_reg_9__5__5_ ( .D(n15183), .CK(clk), .Q(gray_img[1197]) );
  QDFFS gray_img_reg_9__6__5_ ( .D(n15182), .CK(clk), .Q(gray_img[1205]) );
  QDFFS gray_img_reg_9__7__5_ ( .D(n15181), .CK(clk), .Q(gray_img[1213]) );
  QDFFS gray_img_reg_9__8__5_ ( .D(n15180), .CK(clk), .Q(gray_img[1221]) );
  QDFFS gray_img_reg_9__9__5_ ( .D(n15179), .CK(clk), .Q(gray_img[1229]) );
  QDFFS gray_img_reg_9__10__5_ ( .D(n15178), .CK(clk), .Q(gray_img[1237]) );
  QDFFS gray_img_reg_9__11__5_ ( .D(n15177), .CK(clk), .Q(gray_img[1245]) );
  QDFFS gray_img_reg_9__12__5_ ( .D(n15176), .CK(clk), .Q(gray_img[1253]) );
  QDFFS gray_img_reg_9__13__5_ ( .D(n15175), .CK(clk), .Q(gray_img[1261]) );
  QDFFS gray_img_reg_9__14__5_ ( .D(n15174), .CK(clk), .Q(gray_img[1269]) );
  QDFFS gray_img_reg_9__15__5_ ( .D(n15173), .CK(clk), .Q(gray_img[1277]) );
  QDFFS gray_img_reg_10__0__5_ ( .D(n15172), .CK(clk), .Q(gray_img[1285]) );
  QDFFS gray_img_reg_10__1__5_ ( .D(n15171), .CK(clk), .Q(gray_img[1293]) );
  QDFFS gray_img_reg_10__2__5_ ( .D(n15170), .CK(clk), .Q(gray_img[1301]) );
  QDFFS gray_img_reg_10__3__5_ ( .D(n15169), .CK(clk), .Q(gray_img[1309]) );
  QDFFS gray_img_reg_10__4__5_ ( .D(n15168), .CK(clk), .Q(gray_img[1317]) );
  QDFFS gray_img_reg_10__5__5_ ( .D(n15167), .CK(clk), .Q(gray_img[1325]) );
  QDFFS gray_img_reg_10__6__5_ ( .D(n15166), .CK(clk), .Q(gray_img[1333]) );
  QDFFS gray_img_reg_10__7__5_ ( .D(n15165), .CK(clk), .Q(gray_img[1341]) );
  QDFFS gray_img_reg_10__8__5_ ( .D(n15164), .CK(clk), .Q(gray_img[1349]) );
  QDFFS gray_img_reg_10__9__5_ ( .D(n15163), .CK(clk), .Q(gray_img[1357]) );
  QDFFS gray_img_reg_10__10__5_ ( .D(n15162), .CK(clk), .Q(gray_img[1365]) );
  QDFFS gray_img_reg_10__11__5_ ( .D(n15161), .CK(clk), .Q(gray_img[1373]) );
  QDFFS gray_img_reg_10__12__5_ ( .D(n15160), .CK(clk), .Q(gray_img[1381]) );
  QDFFS gray_img_reg_10__13__5_ ( .D(n15159), .CK(clk), .Q(gray_img[1389]) );
  QDFFS gray_img_reg_10__14__5_ ( .D(n15158), .CK(clk), .Q(gray_img[1397]) );
  QDFFS gray_img_reg_10__15__5_ ( .D(n15157), .CK(clk), .Q(gray_img[1405]) );
  QDFFS gray_img_reg_11__0__5_ ( .D(n15156), .CK(clk), .Q(gray_img[1413]) );
  QDFFS gray_img_reg_11__1__5_ ( .D(n15155), .CK(clk), .Q(gray_img[1421]) );
  QDFFS gray_img_reg_11__2__5_ ( .D(n15154), .CK(clk), .Q(gray_img[1429]) );
  QDFFS gray_img_reg_11__3__5_ ( .D(n15153), .CK(clk), .Q(gray_img[1437]) );
  QDFFS gray_img_reg_11__4__5_ ( .D(n15152), .CK(clk), .Q(gray_img[1445]) );
  QDFFS gray_img_reg_11__5__5_ ( .D(n15151), .CK(clk), .Q(gray_img[1453]) );
  QDFFS gray_img_reg_11__6__5_ ( .D(n15150), .CK(clk), .Q(gray_img[1461]) );
  QDFFS gray_img_reg_11__7__5_ ( .D(n15149), .CK(clk), .Q(gray_img[1469]) );
  QDFFS gray_img_reg_11__8__5_ ( .D(n15148), .CK(clk), .Q(gray_img[1477]) );
  QDFFS gray_img_reg_11__9__5_ ( .D(n15147), .CK(clk), .Q(gray_img[1485]) );
  QDFFS gray_img_reg_11__10__5_ ( .D(n15146), .CK(clk), .Q(gray_img[1493]) );
  QDFFS gray_img_reg_11__11__5_ ( .D(n15145), .CK(clk), .Q(gray_img[1501]) );
  QDFFS gray_img_reg_11__12__5_ ( .D(n15144), .CK(clk), .Q(gray_img[1509]) );
  QDFFS gray_img_reg_11__13__5_ ( .D(n15143), .CK(clk), .Q(gray_img[1517]) );
  QDFFS gray_img_reg_11__14__5_ ( .D(n15142), .CK(clk), .Q(gray_img[1525]) );
  QDFFS gray_img_reg_11__15__5_ ( .D(n15141), .CK(clk), .Q(gray_img[1533]) );
  QDFFS gray_img_reg_12__0__5_ ( .D(n15140), .CK(clk), .Q(gray_img[1541]) );
  QDFFS gray_img_reg_12__1__5_ ( .D(n15139), .CK(clk), .Q(gray_img[1549]) );
  QDFFS gray_img_reg_12__2__5_ ( .D(n15138), .CK(clk), .Q(gray_img[1557]) );
  QDFFS gray_img_reg_12__3__5_ ( .D(n15137), .CK(clk), .Q(gray_img[1565]) );
  QDFFS gray_img_reg_12__4__5_ ( .D(n15136), .CK(clk), .Q(gray_img[1573]) );
  QDFFS gray_img_reg_12__5__5_ ( .D(n15135), .CK(clk), .Q(gray_img[1581]) );
  QDFFS gray_img_reg_12__6__5_ ( .D(n15134), .CK(clk), .Q(gray_img[1589]) );
  QDFFS gray_img_reg_12__7__5_ ( .D(n15133), .CK(clk), .Q(gray_img[1597]) );
  QDFFS gray_img_reg_12__8__5_ ( .D(n15132), .CK(clk), .Q(gray_img[1605]) );
  QDFFS gray_img_reg_12__9__5_ ( .D(n15131), .CK(clk), .Q(gray_img[1613]) );
  QDFFS gray_img_reg_12__10__5_ ( .D(n15130), .CK(clk), .Q(gray_img[1621]) );
  QDFFS gray_img_reg_12__11__5_ ( .D(n15129), .CK(clk), .Q(gray_img[1629]) );
  QDFFS gray_img_reg_12__12__5_ ( .D(n15128), .CK(clk), .Q(gray_img[1637]) );
  QDFFS gray_img_reg_12__13__5_ ( .D(n15127), .CK(clk), .Q(gray_img[1645]) );
  QDFFS gray_img_reg_12__14__5_ ( .D(n15126), .CK(clk), .Q(gray_img[1653]) );
  QDFFS gray_img_reg_12__15__5_ ( .D(n15125), .CK(clk), .Q(gray_img[1661]) );
  QDFFS gray_img_reg_13__0__5_ ( .D(n15124), .CK(clk), .Q(gray_img[1669]) );
  QDFFS gray_img_reg_13__1__5_ ( .D(n15123), .CK(clk), .Q(gray_img[1677]) );
  QDFFS gray_img_reg_13__2__5_ ( .D(n15122), .CK(clk), .Q(gray_img[1685]) );
  QDFFS gray_img_reg_13__3__5_ ( .D(n15121), .CK(clk), .Q(gray_img[1693]) );
  QDFFS gray_img_reg_13__4__5_ ( .D(n15120), .CK(clk), .Q(gray_img[1701]) );
  QDFFS gray_img_reg_13__5__5_ ( .D(n15119), .CK(clk), .Q(gray_img[1709]) );
  QDFFS gray_img_reg_13__6__5_ ( .D(n15118), .CK(clk), .Q(gray_img[1717]) );
  QDFFS gray_img_reg_13__7__5_ ( .D(n15117), .CK(clk), .Q(gray_img[1725]) );
  QDFFS gray_img_reg_13__8__5_ ( .D(n15116), .CK(clk), .Q(gray_img[1733]) );
  QDFFS gray_img_reg_13__9__5_ ( .D(n15115), .CK(clk), .Q(gray_img[1741]) );
  QDFFS gray_img_reg_13__10__5_ ( .D(n15114), .CK(clk), .Q(gray_img[1749]) );
  QDFFS gray_img_reg_13__11__5_ ( .D(n15113), .CK(clk), .Q(gray_img[1757]) );
  QDFFS gray_img_reg_13__12__5_ ( .D(n15112), .CK(clk), .Q(gray_img[1765]) );
  QDFFS gray_img_reg_13__13__5_ ( .D(n15111), .CK(clk), .Q(gray_img[1773]) );
  QDFFS gray_img_reg_13__14__5_ ( .D(n15110), .CK(clk), .Q(gray_img[1781]) );
  QDFFS gray_img_reg_13__15__5_ ( .D(n15109), .CK(clk), .Q(gray_img[1789]) );
  QDFFS gray_img_reg_14__0__5_ ( .D(n15108), .CK(clk), .Q(gray_img[1797]) );
  QDFFS gray_img_reg_14__1__5_ ( .D(n15107), .CK(clk), .Q(gray_img[1805]) );
  QDFFS gray_img_reg_14__2__5_ ( .D(n15106), .CK(clk), .Q(gray_img[1813]) );
  QDFFS gray_img_reg_14__3__5_ ( .D(n15105), .CK(clk), .Q(gray_img[1821]) );
  QDFFS gray_img_reg_14__4__5_ ( .D(n15104), .CK(clk), .Q(gray_img[1829]) );
  QDFFS gray_img_reg_14__5__5_ ( .D(n15103), .CK(clk), .Q(gray_img[1837]) );
  QDFFS gray_img_reg_14__6__5_ ( .D(n15102), .CK(clk), .Q(gray_img[1845]) );
  QDFFS gray_img_reg_14__7__5_ ( .D(n15101), .CK(clk), .Q(gray_img[1853]) );
  QDFFS gray_img_reg_14__8__5_ ( .D(n15100), .CK(clk), .Q(gray_img[1861]) );
  QDFFS gray_img_reg_14__9__5_ ( .D(n15099), .CK(clk), .Q(gray_img[1869]) );
  QDFFS gray_img_reg_14__10__5_ ( .D(n15098), .CK(clk), .Q(gray_img[1877]) );
  QDFFS gray_img_reg_14__11__5_ ( .D(n15097), .CK(clk), .Q(gray_img[1885]) );
  QDFFS gray_img_reg_14__12__5_ ( .D(n15096), .CK(clk), .Q(gray_img[1893]) );
  QDFFS gray_img_reg_14__13__5_ ( .D(n15095), .CK(clk), .Q(gray_img[1901]) );
  QDFFS gray_img_reg_14__14__5_ ( .D(n15094), .CK(clk), .Q(gray_img[1909]) );
  QDFFS gray_img_reg_14__15__5_ ( .D(n15093), .CK(clk), .Q(gray_img[1917]) );
  QDFFS gray_img_reg_15__0__5_ ( .D(n15092), .CK(clk), .Q(gray_img[1925]) );
  QDFFS gray_img_reg_15__1__5_ ( .D(n15091), .CK(clk), .Q(gray_img[1933]) );
  QDFFS gray_img_reg_15__2__5_ ( .D(n15090), .CK(clk), .Q(gray_img[1941]) );
  QDFFS gray_img_reg_15__3__5_ ( .D(n15089), .CK(clk), .Q(gray_img[1949]) );
  QDFFS gray_img_reg_15__4__5_ ( .D(n15088), .CK(clk), .Q(gray_img[1957]) );
  QDFFS gray_img_reg_15__5__5_ ( .D(n15087), .CK(clk), .Q(gray_img[1965]) );
  QDFFS gray_img_reg_15__6__5_ ( .D(n15086), .CK(clk), .Q(gray_img[1973]) );
  QDFFS gray_img_reg_15__7__5_ ( .D(n15085), .CK(clk), .Q(gray_img[1981]) );
  QDFFS gray_img_reg_15__8__5_ ( .D(n15084), .CK(clk), .Q(gray_img[1989]) );
  QDFFS gray_img_reg_15__9__5_ ( .D(n15083), .CK(clk), .Q(gray_img[1997]) );
  QDFFS gray_img_reg_15__10__5_ ( .D(n15082), .CK(clk), .Q(gray_img[2005]) );
  QDFFS gray_img_reg_15__11__5_ ( .D(n15081), .CK(clk), .Q(gray_img[2013]) );
  QDFFS gray_img_reg_15__12__5_ ( .D(n15080), .CK(clk), .Q(gray_img[2021]) );
  QDFFS gray_img_reg_15__13__5_ ( .D(n15079), .CK(clk), .Q(gray_img[2029]) );
  QDFFS gray_img_reg_15__14__5_ ( .D(n15078), .CK(clk), .Q(gray_img[2037]) );
  QDFFS gray_img_reg_15__15__5_ ( .D(n15077), .CK(clk), .Q(gray_img[2045]) );
  QDFFS gray_img_reg_7__3__5_ ( .D(n15073), .CK(clk), .Q(gray_img[925]) );
  QDFFS gray_img_reg_0__4__5_ ( .D(n14252), .CK(clk), .Q(gray_img[37]) );
  QDFFS gray_img_reg_0__5__5_ ( .D(n14243), .CK(clk), .Q(gray_img[45]) );
  QDFFS gray_img_reg_0__6__5_ ( .D(n14234), .CK(clk), .Q(gray_img[53]) );
  QDFFS gray_img_reg_0__7__5_ ( .D(n14225), .CK(clk), .Q(gray_img[61]) );
  QDFFS gray_img_reg_1__4__5_ ( .D(n14208), .CK(clk), .Q(gray_img[165]) );
  QDFFS gray_img_reg_1__5__5_ ( .D(n14199), .CK(clk), .Q(gray_img[173]) );
  QDFFS gray_img_reg_1__6__5_ ( .D(n14190), .CK(clk), .Q(gray_img[181]) );
  QDFFS gray_img_reg_1__7__5_ ( .D(n14181), .CK(clk), .Q(gray_img[189]) );
  QDFFS gray_img_reg_2__4__5_ ( .D(n14164), .CK(clk), .Q(gray_img[293]) );
  QDFFS gray_img_reg_2__5__5_ ( .D(n14155), .CK(clk), .Q(gray_img[301]) );
  QDFFS gray_img_reg_2__6__5_ ( .D(n14146), .CK(clk), .Q(gray_img[309]) );
  QDFFS gray_img_reg_2__7__5_ ( .D(n14137), .CK(clk), .Q(gray_img[317]) );
  QDFFS gray_img_reg_3__4__5_ ( .D(n14120), .CK(clk), .Q(gray_img[421]) );
  QDFFS gray_img_reg_3__5__5_ ( .D(n14111), .CK(clk), .Q(gray_img[429]) );
  QDFFS gray_img_reg_3__6__5_ ( .D(n14102), .CK(clk), .Q(gray_img[437]) );
  QDFFS gray_img_reg_3__7__5_ ( .D(n14093), .CK(clk), .Q(gray_img[445]) );
  QDFFS gray_img_reg_4__0__5_ ( .D(n14068), .CK(clk), .Q(gray_img[517]) );
  QDFFS gray_img_reg_4__1__5_ ( .D(n14059), .CK(clk), .Q(gray_img[525]) );
  QDFFS gray_img_reg_4__2__5_ ( .D(n14050), .CK(clk), .Q(gray_img[533]) );
  QDFFS gray_img_reg_4__3__5_ ( .D(n14041), .CK(clk), .Q(gray_img[541]) );
  QDFFS gray_img_reg_4__4__5_ ( .D(n14032), .CK(clk), .Q(gray_img[549]) );
  QDFFS gray_img_reg_4__5__5_ ( .D(n14023), .CK(clk), .Q(gray_img[557]) );
  QDFFS gray_img_reg_4__6__5_ ( .D(n14014), .CK(clk), .Q(gray_img[565]) );
  QDFFS gray_img_reg_4__7__5_ ( .D(n14005), .CK(clk), .Q(gray_img[573]) );
  QDFFS gray_img_reg_5__0__5_ ( .D(n13980), .CK(clk), .Q(gray_img[645]) );
  QDFFS gray_img_reg_5__1__5_ ( .D(n13971), .CK(clk), .Q(gray_img[653]) );
  QDFFS gray_img_reg_5__2__5_ ( .D(n13962), .CK(clk), .Q(gray_img[661]) );
  QDFFS gray_img_reg_5__3__5_ ( .D(n13954), .CK(clk), .Q(gray_img[669]) );
  QDFFS gray_img_reg_5__4__5_ ( .D(n13946), .CK(clk), .Q(gray_img[677]) );
  QDFFS gray_img_reg_5__5__5_ ( .D(n13939), .CK(clk), .Q(gray_img[685]) );
  QDFFS gray_img_reg_5__6__5_ ( .D(n13932), .CK(clk), .Q(gray_img[693]) );
  QDFFS gray_img_reg_5__7__5_ ( .D(n13926), .CK(clk), .Q(gray_img[701]) );
  QDFFS gray_img_reg_6__0__5_ ( .D(n13904), .CK(clk), .Q(gray_img[773]) );
  QDFFS gray_img_reg_6__1__5_ ( .D(n13898), .CK(clk), .Q(gray_img[781]) );
  QDFFS gray_img_reg_6__2__5_ ( .D(n13892), .CK(clk), .Q(gray_img[789]) );
  QDFFS gray_img_reg_6__3__5_ ( .D(n13886), .CK(clk), .Q(gray_img[797]) );
  QDFFS gray_img_reg_6__4__5_ ( .D(n13880), .CK(clk), .Q(gray_img[805]) );
  QDFFS gray_img_reg_6__5__5_ ( .D(n13874), .CK(clk), .Q(gray_img[813]) );
  QDFFS gray_img_reg_6__6__5_ ( .D(n13868), .CK(clk), .Q(gray_img[821]) );
  QDFFS gray_img_reg_6__7__5_ ( .D(n13862), .CK(clk), .Q(gray_img[829]) );
  QDFFS gray_img_reg_7__0__5_ ( .D(n13840), .CK(clk), .Q(gray_img[901]) );
  QDFFS gray_img_reg_7__1__5_ ( .D(n13835), .CK(clk), .Q(gray_img[909]) );
  QDFFS gray_img_reg_7__2__5_ ( .D(n13830), .CK(clk), .Q(gray_img[917]) );
  QDFFS gray_img_reg_3__1__5_ ( .D(n15072), .CK(clk), .Q(gray_img[397]) );
  QDFFS gray_img_reg_0__2__5_ ( .D(n13797), .CK(clk), .Q(gray_img[21]) );
  QDFFS gray_img_reg_0__3__5_ ( .D(n13787), .CK(clk), .Q(gray_img[29]) );
  QDFFS gray_img_reg_1__2__5_ ( .D(n13767), .CK(clk), .Q(gray_img[149]) );
  QDFFS gray_img_reg_1__3__5_ ( .D(n13757), .CK(clk), .Q(gray_img[157]) );
  QDFFS gray_img_reg_0__1__5_ ( .D(n13749), .CK(clk), .Q(gray_img[13]) );
  QDFFS gray_img_reg_2__0__5_ ( .D(n13731), .CK(clk), .Q(gray_img[261]) );
  QDFFS gray_img_reg_2__1__5_ ( .D(n13702), .CK(clk), .Q(gray_img[269]) );
  QDFFS gray_img_reg_2__2__5_ ( .D(n13676), .CK(clk), .Q(gray_img[277]) );
  QDFFS gray_img_reg_2__3__5_ ( .D(n13653), .CK(clk), .Q(gray_img[285]) );
  QDFFS gray_img_reg_3__0__5_ ( .D(n13633), .CK(clk), .Q(gray_img[389]) );
  QDFFS gray_img_reg_1__0__5_ ( .D(n13624), .CK(clk), .Q(gray_img[133]) );
  QDFFS gray_img_reg_7__4__5_ ( .D(n13621), .CK(clk), .Q(gray_img[933]) );
  QDFFS gray_img_reg_7__5__5_ ( .D(n13620), .CK(clk), .Q(gray_img[941]) );
  QDFFS gray_img_reg_3__2__5_ ( .D(n15269), .CK(clk), .Q(gray_img[405]) );
  QDFFS gray_img_reg_7__6__5_ ( .D(n13619), .CK(clk), .Q(gray_img[949]) );
  QDFFS gray_img_reg_7__7__5_ ( .D(n13618), .CK(clk), .Q(gray_img[957]) );
  QDFFS gray_img_reg_3__3__5_ ( .D(n15074), .CK(clk), .Q(gray_img[413]) );
  QDFFS gray_img_reg_1__1__5_ ( .D(n15075), .CK(clk), .Q(gray_img[141]) );
  QDFFS gray_img_reg_0__0__4_ ( .D(n14876), .CK(clk), .Q(gray_img[4]) );
  QDFFS mem_data_out_reg_shift_0_reg_0__4_ ( .D(n15811), .CK(clk), .Q(
        mem_data_out_reg_shift_0[4]) );
  QDFFS mem_data_out_reg_shift_0_reg_1__4_ ( .D(mem_data_out_reg_shift_0[4]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[12]) );
  QDFFS mem_data_out_reg_shift_0_reg_2__4_ ( .D(mem_data_out_reg_shift_0[12]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[20]) );
  QDFFS mem_data_out_reg_shift_0_reg_3__4_ ( .D(mem_data_out_reg_shift_0[20]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[28]) );
  QDFFS mem_data_out_reg_shift_0_reg_4__4_ ( .D(mem_data_out_reg_shift_0[28]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[36]) );
  QDFFS mem_data_out_reg_shift_0_reg_5__4_ ( .D(mem_data_out_reg_shift_0[36]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[44]) );
  QDFFS mem_data_out_reg_shift_0_reg_6__4_ ( .D(mem_data_out_reg_shift_0[44]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[52]) );
  QDFFS mem_data_out_reg_shift_0_reg_7__4_ ( .D(mem_data_out_reg_shift_0[52]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[60]) );
  QDFFS mem_data_out_reg_shift_0_reg_8__4_ ( .D(mem_data_out_reg_shift_0[60]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[68]) );
  QDFFS mem_data_out_reg_shift_0_reg_9__4_ ( .D(mem_data_out_reg_shift_0[68]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[76]) );
  QDFFS mem_data_out_reg_shift_0_reg_10__4_ ( .D(mem_data_out_reg_shift_0[76]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[84]) );
  QDFFS mem_data_out_reg_shift_0_reg_11__4_ ( .D(mem_data_out_reg_shift_0[84]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[92]) );
  QDFFS mem_data_out_reg_shift_0_reg_12__4_ ( .D(mem_data_out_reg_shift_0[92]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[100]) );
  QDFFS mem_data_out_reg_shift_0_reg_13__4_ ( .D(mem_data_out_reg_shift_0[100]), .CK(clk), .Q(mem_data_out_reg_shift_0[108]) );
  QDFFS mem_data_out_reg_shift_0_reg_14__4_ ( .D(mem_data_out_reg_shift_0[108]), .CK(clk), .Q(mem_data_out_reg_shift_0[116]) );
  QDFFS mem_data_out_reg_shift_0_reg_15__4_ ( .D(mem_data_out_reg_shift_0[116]), .CK(clk), .Q(mem_data_out_reg_shift_0[124]) );
  QDFFS mem_data_out_reg_shift_1_reg_0__4_ ( .D(n15828), .CK(clk), .Q(
        mem_data_out_reg_shift_1[4]) );
  QDFFS mem_data_out_reg_shift_1_reg_1__4_ ( .D(mem_data_out_reg_shift_1[4]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[12]) );
  QDFFS mem_data_out_reg_shift_1_reg_3__4_ ( .D(mem_data_out_reg_shift_1[20]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[28]) );
  QDFFS mem_data_out_reg_shift_1_reg_4__4_ ( .D(mem_data_out_reg_shift_1[28]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[36]) );
  QDFFS mem_data_out_reg_shift_1_reg_5__4_ ( .D(mem_data_out_reg_shift_1[36]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[44]) );
  QDFFS mem_data_out_reg_shift_1_reg_6__4_ ( .D(mem_data_out_reg_shift_1[44]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[52]) );
  QDFFS mem_data_out_reg_shift_1_reg_7__4_ ( .D(mem_data_out_reg_shift_1[52]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[60]) );
  QDFFS mem_data_out_reg_shift_1_reg_8__4_ ( .D(mem_data_out_reg_shift_1[60]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[68]) );
  QDFFS mem_data_out_reg_shift_1_reg_9__4_ ( .D(mem_data_out_reg_shift_1[68]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[76]) );
  QDFFS mem_data_out_reg_shift_1_reg_10__4_ ( .D(mem_data_out_reg_shift_1[76]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[84]) );
  QDFFS mem_data_out_reg_shift_1_reg_11__4_ ( .D(mem_data_out_reg_shift_1[84]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[92]) );
  QDFFS mem_data_out_reg_shift_1_reg_12__4_ ( .D(mem_data_out_reg_shift_1[92]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[100]) );
  QDFFS mem_data_out_reg_shift_1_reg_13__4_ ( .D(mem_data_out_reg_shift_1[100]), .CK(clk), .Q(mem_data_out_reg_shift_1[108]) );
  QDFFS mem_data_out_reg_shift_1_reg_14__4_ ( .D(mem_data_out_reg_shift_1[108]), .CK(clk), .Q(mem_data_out_reg_shift_1[116]) );
  QDFFS mem_data_out_reg_shift_1_reg_15__4_ ( .D(mem_data_out_reg_shift_1[116]), .CK(clk), .Q(mem_data_out_reg_shift_1[124]) );
  QDFFS mem_data_out_reg_shift_2_reg_0__4_ ( .D(n15836), .CK(clk), .Q(
        mem_data_out_reg_shift_2[4]) );
  QDFFS mem_data_out_reg_shift_2_reg_1__4_ ( .D(mem_data_out_reg_shift_2[4]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[12]) );
  QDFFS mem_data_out_reg_shift_2_reg_2__4_ ( .D(mem_data_out_reg_shift_2[12]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[20]) );
  QDFFS mem_data_out_reg_shift_2_reg_3__4_ ( .D(mem_data_out_reg_shift_2[20]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[28]) );
  QDFFS gray_img_reg_0__8__4_ ( .D(n15068), .CK(clk), .Q(gray_img[68]) );
  QDFFS gray_img_reg_0__9__4_ ( .D(n15067), .CK(clk), .Q(gray_img[76]) );
  QDFFS gray_img_reg_0__10__4_ ( .D(n15066), .CK(clk), .Q(gray_img[84]) );
  QDFFS gray_img_reg_0__11__4_ ( .D(n15065), .CK(clk), .Q(gray_img[92]) );
  QDFFS gray_img_reg_0__12__4_ ( .D(n15064), .CK(clk), .Q(gray_img[100]) );
  QDFFS gray_img_reg_0__13__4_ ( .D(n15063), .CK(clk), .Q(gray_img[108]) );
  QDFFS gray_img_reg_0__14__4_ ( .D(n15062), .CK(clk), .Q(gray_img[116]) );
  QDFFS gray_img_reg_0__15__4_ ( .D(n15061), .CK(clk), .Q(gray_img[124]) );
  QDFFS gray_img_reg_1__8__4_ ( .D(n15060), .CK(clk), .Q(gray_img[196]) );
  QDFFS gray_img_reg_1__9__4_ ( .D(n15059), .CK(clk), .Q(gray_img[204]) );
  QDFFS gray_img_reg_1__10__4_ ( .D(n15058), .CK(clk), .Q(gray_img[212]) );
  QDFFS gray_img_reg_1__11__4_ ( .D(n15057), .CK(clk), .Q(gray_img[220]) );
  QDFFS gray_img_reg_1__12__4_ ( .D(n15056), .CK(clk), .Q(gray_img[228]) );
  QDFFS gray_img_reg_1__13__4_ ( .D(n15055), .CK(clk), .Q(gray_img[236]) );
  QDFFS gray_img_reg_1__14__4_ ( .D(n15054), .CK(clk), .Q(gray_img[244]) );
  QDFFS gray_img_reg_1__15__4_ ( .D(n15053), .CK(clk), .Q(gray_img[252]) );
  QDFFS gray_img_reg_2__8__4_ ( .D(n15052), .CK(clk), .Q(gray_img[324]) );
  QDFFS gray_img_reg_2__9__4_ ( .D(n15051), .CK(clk), .Q(gray_img[332]) );
  QDFFS gray_img_reg_2__10__4_ ( .D(n15050), .CK(clk), .Q(gray_img[340]) );
  QDFFS gray_img_reg_2__11__4_ ( .D(n15049), .CK(clk), .Q(gray_img[348]) );
  QDFFS gray_img_reg_2__12__4_ ( .D(n15048), .CK(clk), .Q(gray_img[356]) );
  QDFFS gray_img_reg_2__13__4_ ( .D(n15047), .CK(clk), .Q(gray_img[364]) );
  QDFFS gray_img_reg_2__14__4_ ( .D(n15046), .CK(clk), .Q(gray_img[372]) );
  QDFFS gray_img_reg_2__15__4_ ( .D(n15045), .CK(clk), .Q(gray_img[380]) );
  QDFFS gray_img_reg_3__8__4_ ( .D(n15044), .CK(clk), .Q(gray_img[452]) );
  QDFFS gray_img_reg_3__9__4_ ( .D(n15043), .CK(clk), .Q(gray_img[460]) );
  QDFFS gray_img_reg_3__10__4_ ( .D(n15042), .CK(clk), .Q(gray_img[468]) );
  QDFFS gray_img_reg_3__11__4_ ( .D(n15041), .CK(clk), .Q(gray_img[476]) );
  QDFFS gray_img_reg_3__12__4_ ( .D(n15040), .CK(clk), .Q(gray_img[484]) );
  QDFFS gray_img_reg_3__13__4_ ( .D(n15039), .CK(clk), .Q(gray_img[492]) );
  QDFFS gray_img_reg_3__14__4_ ( .D(n15038), .CK(clk), .Q(gray_img[500]) );
  QDFFS gray_img_reg_3__15__4_ ( .D(n15037), .CK(clk), .Q(gray_img[508]) );
  QDFFS gray_img_reg_4__8__4_ ( .D(n15036), .CK(clk), .Q(gray_img[580]) );
  QDFFS gray_img_reg_4__9__4_ ( .D(n15035), .CK(clk), .Q(gray_img[588]) );
  QDFFS gray_img_reg_4__10__4_ ( .D(n15034), .CK(clk), .Q(gray_img[596]) );
  QDFFS gray_img_reg_4__11__4_ ( .D(n15033), .CK(clk), .Q(gray_img[604]) );
  QDFFS gray_img_reg_4__12__4_ ( .D(n15032), .CK(clk), .Q(gray_img[612]) );
  QDFFS gray_img_reg_4__13__4_ ( .D(n15031), .CK(clk), .Q(gray_img[620]) );
  QDFFS gray_img_reg_4__14__4_ ( .D(n15030), .CK(clk), .Q(gray_img[628]) );
  QDFFS gray_img_reg_4__15__4_ ( .D(n15029), .CK(clk), .Q(gray_img[636]) );
  QDFFS gray_img_reg_5__8__4_ ( .D(n15028), .CK(clk), .Q(gray_img[708]) );
  QDFFS gray_img_reg_5__9__4_ ( .D(n15027), .CK(clk), .Q(gray_img[716]) );
  QDFFS gray_img_reg_5__10__4_ ( .D(n15026), .CK(clk), .Q(gray_img[724]) );
  QDFFS gray_img_reg_5__11__4_ ( .D(n15025), .CK(clk), .Q(gray_img[732]) );
  QDFFS gray_img_reg_5__12__4_ ( .D(n15024), .CK(clk), .Q(gray_img[740]) );
  QDFFS gray_img_reg_5__13__4_ ( .D(n15023), .CK(clk), .Q(gray_img[748]) );
  QDFFS gray_img_reg_5__14__4_ ( .D(n15022), .CK(clk), .Q(gray_img[756]) );
  QDFFS gray_img_reg_5__15__4_ ( .D(n15021), .CK(clk), .Q(gray_img[764]) );
  QDFFS gray_img_reg_6__8__4_ ( .D(n15020), .CK(clk), .Q(gray_img[836]) );
  QDFFS gray_img_reg_6__9__4_ ( .D(n15019), .CK(clk), .Q(gray_img[844]) );
  QDFFS gray_img_reg_6__10__4_ ( .D(n15018), .CK(clk), .Q(gray_img[852]) );
  QDFFS gray_img_reg_6__11__4_ ( .D(n15017), .CK(clk), .Q(gray_img[860]) );
  QDFFS gray_img_reg_6__12__4_ ( .D(n15016), .CK(clk), .Q(gray_img[868]) );
  QDFFS gray_img_reg_6__13__4_ ( .D(n15015), .CK(clk), .Q(gray_img[876]) );
  QDFFS gray_img_reg_6__14__4_ ( .D(n15014), .CK(clk), .Q(gray_img[884]) );
  QDFFS gray_img_reg_6__15__4_ ( .D(n15013), .CK(clk), .Q(gray_img[892]) );
  QDFFS gray_img_reg_7__8__4_ ( .D(n15012), .CK(clk), .Q(gray_img[964]) );
  QDFFS gray_img_reg_7__9__4_ ( .D(n15011), .CK(clk), .Q(gray_img[972]) );
  QDFFS gray_img_reg_7__10__4_ ( .D(n15010), .CK(clk), .Q(gray_img[980]) );
  QDFFS gray_img_reg_7__11__4_ ( .D(n15009), .CK(clk), .Q(gray_img[988]) );
  QDFFS gray_img_reg_7__12__4_ ( .D(n15008), .CK(clk), .Q(gray_img[996]) );
  QDFFS gray_img_reg_7__13__4_ ( .D(n15007), .CK(clk), .Q(gray_img[1004]) );
  QDFFS gray_img_reg_7__14__4_ ( .D(n15006), .CK(clk), .Q(gray_img[1012]) );
  QDFFS gray_img_reg_7__15__4_ ( .D(n15005), .CK(clk), .Q(gray_img[1020]) );
  QDFFS gray_img_reg_8__0__4_ ( .D(n15004), .CK(clk), .Q(gray_img[1028]) );
  QDFFS gray_img_reg_8__1__4_ ( .D(n15003), .CK(clk), .Q(gray_img[1036]) );
  QDFFS gray_img_reg_8__2__4_ ( .D(n15002), .CK(clk), .Q(gray_img[1044]) );
  QDFFS gray_img_reg_8__3__4_ ( .D(n15001), .CK(clk), .Q(gray_img[1052]) );
  QDFFS gray_img_reg_8__4__4_ ( .D(n15000), .CK(clk), .Q(gray_img[1060]) );
  QDFFS gray_img_reg_8__5__4_ ( .D(n14999), .CK(clk), .Q(gray_img[1068]) );
  QDFFS gray_img_reg_8__6__4_ ( .D(n14998), .CK(clk), .Q(gray_img[1076]) );
  QDFFS gray_img_reg_8__7__4_ ( .D(n14997), .CK(clk), .Q(gray_img[1084]) );
  QDFFS gray_img_reg_8__8__4_ ( .D(n14996), .CK(clk), .Q(gray_img[1092]) );
  QDFFS gray_img_reg_8__9__4_ ( .D(n14995), .CK(clk), .Q(gray_img[1100]) );
  QDFFS gray_img_reg_8__10__4_ ( .D(n14994), .CK(clk), .Q(gray_img[1108]) );
  QDFFS gray_img_reg_8__11__4_ ( .D(n14993), .CK(clk), .Q(gray_img[1116]) );
  QDFFS gray_img_reg_8__12__4_ ( .D(n14992), .CK(clk), .Q(gray_img[1124]) );
  QDFFS gray_img_reg_8__13__4_ ( .D(n14991), .CK(clk), .Q(gray_img[1132]) );
  QDFFS gray_img_reg_8__14__4_ ( .D(n14990), .CK(clk), .Q(gray_img[1140]) );
  QDFFS gray_img_reg_8__15__4_ ( .D(n14989), .CK(clk), .Q(gray_img[1148]) );
  QDFFS gray_img_reg_9__0__4_ ( .D(n14988), .CK(clk), .Q(gray_img[1156]) );
  QDFFS gray_img_reg_9__1__4_ ( .D(n14987), .CK(clk), .Q(gray_img[1164]) );
  QDFFS gray_img_reg_9__2__4_ ( .D(n14986), .CK(clk), .Q(gray_img[1172]) );
  QDFFS gray_img_reg_9__3__4_ ( .D(n14985), .CK(clk), .Q(gray_img[1180]) );
  QDFFS gray_img_reg_9__4__4_ ( .D(n14984), .CK(clk), .Q(gray_img[1188]) );
  QDFFS gray_img_reg_9__5__4_ ( .D(n14983), .CK(clk), .Q(gray_img[1196]) );
  QDFFS gray_img_reg_9__6__4_ ( .D(n14982), .CK(clk), .Q(gray_img[1204]) );
  QDFFS gray_img_reg_9__7__4_ ( .D(n14981), .CK(clk), .Q(gray_img[1212]) );
  QDFFS gray_img_reg_9__8__4_ ( .D(n14980), .CK(clk), .Q(gray_img[1220]) );
  QDFFS gray_img_reg_9__9__4_ ( .D(n14979), .CK(clk), .Q(gray_img[1228]) );
  QDFFS gray_img_reg_9__10__4_ ( .D(n14978), .CK(clk), .Q(gray_img[1236]) );
  QDFFS gray_img_reg_9__11__4_ ( .D(n14977), .CK(clk), .Q(gray_img[1244]) );
  QDFFS gray_img_reg_9__12__4_ ( .D(n14976), .CK(clk), .Q(gray_img[1252]) );
  QDFFS gray_img_reg_9__13__4_ ( .D(n14975), .CK(clk), .Q(gray_img[1260]) );
  QDFFS gray_img_reg_9__14__4_ ( .D(n14974), .CK(clk), .Q(gray_img[1268]) );
  QDFFS gray_img_reg_9__15__4_ ( .D(n14973), .CK(clk), .Q(gray_img[1276]) );
  QDFFS gray_img_reg_10__0__4_ ( .D(n14972), .CK(clk), .Q(gray_img[1284]) );
  QDFFS gray_img_reg_10__1__4_ ( .D(n14971), .CK(clk), .Q(gray_img[1292]) );
  QDFFS gray_img_reg_10__2__4_ ( .D(n14970), .CK(clk), .Q(gray_img[1300]) );
  QDFFS gray_img_reg_10__3__4_ ( .D(n14969), .CK(clk), .Q(gray_img[1308]) );
  QDFFS gray_img_reg_10__4__4_ ( .D(n14968), .CK(clk), .Q(gray_img[1316]) );
  QDFFS gray_img_reg_10__5__4_ ( .D(n14967), .CK(clk), .Q(gray_img[1324]) );
  QDFFS gray_img_reg_10__6__4_ ( .D(n14966), .CK(clk), .Q(gray_img[1332]) );
  QDFFS gray_img_reg_10__7__4_ ( .D(n14965), .CK(clk), .Q(gray_img[1340]) );
  QDFFS gray_img_reg_10__8__4_ ( .D(n14964), .CK(clk), .Q(gray_img[1348]) );
  QDFFS gray_img_reg_10__9__4_ ( .D(n14963), .CK(clk), .Q(gray_img[1356]) );
  QDFFS gray_img_reg_10__10__4_ ( .D(n14962), .CK(clk), .Q(gray_img[1364]) );
  QDFFS gray_img_reg_10__11__4_ ( .D(n14961), .CK(clk), .Q(gray_img[1372]) );
  QDFFS gray_img_reg_10__12__4_ ( .D(n14960), .CK(clk), .Q(gray_img[1380]) );
  QDFFS gray_img_reg_10__13__4_ ( .D(n14959), .CK(clk), .Q(gray_img[1388]) );
  QDFFS gray_img_reg_10__14__4_ ( .D(n14958), .CK(clk), .Q(gray_img[1396]) );
  QDFFS gray_img_reg_10__15__4_ ( .D(n14957), .CK(clk), .Q(gray_img[1404]) );
  QDFFS gray_img_reg_11__0__4_ ( .D(n14956), .CK(clk), .Q(gray_img[1412]) );
  QDFFS gray_img_reg_11__1__4_ ( .D(n14955), .CK(clk), .Q(gray_img[1420]) );
  QDFFS gray_img_reg_11__2__4_ ( .D(n14954), .CK(clk), .Q(gray_img[1428]) );
  QDFFS gray_img_reg_11__3__4_ ( .D(n14953), .CK(clk), .Q(gray_img[1436]) );
  QDFFS gray_img_reg_11__4__4_ ( .D(n14952), .CK(clk), .Q(gray_img[1444]) );
  QDFFS gray_img_reg_11__5__4_ ( .D(n14951), .CK(clk), .Q(gray_img[1452]) );
  QDFFS gray_img_reg_11__6__4_ ( .D(n14950), .CK(clk), .Q(gray_img[1460]) );
  QDFFS gray_img_reg_11__7__4_ ( .D(n14949), .CK(clk), .Q(gray_img[1468]) );
  QDFFS gray_img_reg_11__8__4_ ( .D(n14948), .CK(clk), .Q(gray_img[1476]) );
  QDFFS gray_img_reg_11__9__4_ ( .D(n14947), .CK(clk), .Q(gray_img[1484]) );
  QDFFS gray_img_reg_11__10__4_ ( .D(n14946), .CK(clk), .Q(gray_img[1492]) );
  QDFFS gray_img_reg_11__11__4_ ( .D(n14945), .CK(clk), .Q(gray_img[1500]) );
  QDFFS gray_img_reg_11__12__4_ ( .D(n14944), .CK(clk), .Q(gray_img[1508]) );
  QDFFS gray_img_reg_11__13__4_ ( .D(n14943), .CK(clk), .Q(gray_img[1516]) );
  QDFFS gray_img_reg_11__14__4_ ( .D(n14942), .CK(clk), .Q(gray_img[1524]) );
  QDFFS gray_img_reg_11__15__4_ ( .D(n14941), .CK(clk), .Q(gray_img[1532]) );
  QDFFS gray_img_reg_12__0__4_ ( .D(n14940), .CK(clk), .Q(gray_img[1540]) );
  QDFFS gray_img_reg_12__1__4_ ( .D(n14939), .CK(clk), .Q(gray_img[1548]) );
  QDFFS gray_img_reg_12__2__4_ ( .D(n14938), .CK(clk), .Q(gray_img[1556]) );
  QDFFS gray_img_reg_12__3__4_ ( .D(n14937), .CK(clk), .Q(gray_img[1564]) );
  QDFFS gray_img_reg_12__4__4_ ( .D(n14936), .CK(clk), .Q(gray_img[1572]) );
  QDFFS gray_img_reg_12__5__4_ ( .D(n14935), .CK(clk), .Q(gray_img[1580]) );
  QDFFS gray_img_reg_12__6__4_ ( .D(n14934), .CK(clk), .Q(gray_img[1588]) );
  QDFFS gray_img_reg_12__7__4_ ( .D(n14933), .CK(clk), .Q(gray_img[1596]) );
  QDFFS gray_img_reg_12__8__4_ ( .D(n14932), .CK(clk), .Q(gray_img[1604]) );
  QDFFS gray_img_reg_12__9__4_ ( .D(n14931), .CK(clk), .Q(gray_img[1612]) );
  QDFFS gray_img_reg_12__10__4_ ( .D(n14930), .CK(clk), .Q(gray_img[1620]) );
  QDFFS gray_img_reg_12__11__4_ ( .D(n14929), .CK(clk), .Q(gray_img[1628]) );
  QDFFS gray_img_reg_12__12__4_ ( .D(n14928), .CK(clk), .Q(gray_img[1636]) );
  QDFFS gray_img_reg_12__13__4_ ( .D(n14927), .CK(clk), .Q(gray_img[1644]) );
  QDFFS gray_img_reg_12__14__4_ ( .D(n14926), .CK(clk), .Q(gray_img[1652]) );
  QDFFS gray_img_reg_12__15__4_ ( .D(n14925), .CK(clk), .Q(gray_img[1660]) );
  QDFFS gray_img_reg_13__0__4_ ( .D(n14924), .CK(clk), .Q(gray_img[1668]) );
  QDFFS gray_img_reg_13__1__4_ ( .D(n14923), .CK(clk), .Q(gray_img[1676]) );
  QDFFS gray_img_reg_13__2__4_ ( .D(n14922), .CK(clk), .Q(gray_img[1684]) );
  QDFFS gray_img_reg_13__3__4_ ( .D(n14921), .CK(clk), .Q(gray_img[1692]) );
  QDFFS gray_img_reg_13__4__4_ ( .D(n14920), .CK(clk), .Q(gray_img[1700]) );
  QDFFS gray_img_reg_13__5__4_ ( .D(n14919), .CK(clk), .Q(gray_img[1708]) );
  QDFFS gray_img_reg_13__6__4_ ( .D(n14918), .CK(clk), .Q(gray_img[1716]) );
  QDFFS gray_img_reg_13__7__4_ ( .D(n14917), .CK(clk), .Q(gray_img[1724]) );
  QDFFS gray_img_reg_13__8__4_ ( .D(n14916), .CK(clk), .Q(gray_img[1732]) );
  QDFFS gray_img_reg_13__9__4_ ( .D(n14915), .CK(clk), .Q(gray_img[1740]) );
  QDFFS gray_img_reg_13__10__4_ ( .D(n14914), .CK(clk), .Q(gray_img[1748]) );
  QDFFS gray_img_reg_13__11__4_ ( .D(n14913), .CK(clk), .Q(gray_img[1756]) );
  QDFFS gray_img_reg_13__12__4_ ( .D(n14912), .CK(clk), .Q(gray_img[1764]) );
  QDFFS gray_img_reg_13__13__4_ ( .D(n14911), .CK(clk), .Q(gray_img[1772]) );
  QDFFS gray_img_reg_13__14__4_ ( .D(n14910), .CK(clk), .Q(gray_img[1780]) );
  QDFFS gray_img_reg_13__15__4_ ( .D(n14909), .CK(clk), .Q(gray_img[1788]) );
  QDFFS gray_img_reg_14__0__4_ ( .D(n14908), .CK(clk), .Q(gray_img[1796]) );
  QDFFS gray_img_reg_14__1__4_ ( .D(n14907), .CK(clk), .Q(gray_img[1804]) );
  QDFFS gray_img_reg_14__2__4_ ( .D(n14906), .CK(clk), .Q(gray_img[1812]) );
  QDFFS gray_img_reg_14__3__4_ ( .D(n14905), .CK(clk), .Q(gray_img[1820]) );
  QDFFS gray_img_reg_14__4__4_ ( .D(n14904), .CK(clk), .Q(gray_img[1828]) );
  QDFFS gray_img_reg_14__5__4_ ( .D(n14903), .CK(clk), .Q(gray_img[1836]) );
  QDFFS gray_img_reg_14__6__4_ ( .D(n14902), .CK(clk), .Q(gray_img[1844]) );
  QDFFS gray_img_reg_14__7__4_ ( .D(n14901), .CK(clk), .Q(gray_img[1852]) );
  QDFFS gray_img_reg_14__8__4_ ( .D(n14900), .CK(clk), .Q(gray_img[1860]) );
  QDFFS gray_img_reg_14__9__4_ ( .D(n14899), .CK(clk), .Q(gray_img[1868]) );
  QDFFS gray_img_reg_14__10__4_ ( .D(n14898), .CK(clk), .Q(gray_img[1876]) );
  QDFFS gray_img_reg_14__11__4_ ( .D(n14897), .CK(clk), .Q(gray_img[1884]) );
  QDFFS gray_img_reg_14__12__4_ ( .D(n14896), .CK(clk), .Q(gray_img[1892]) );
  QDFFS gray_img_reg_14__13__4_ ( .D(n14895), .CK(clk), .Q(gray_img[1900]) );
  QDFFS gray_img_reg_14__14__4_ ( .D(n14894), .CK(clk), .Q(gray_img[1908]) );
  QDFFS gray_img_reg_14__15__4_ ( .D(n14893), .CK(clk), .Q(gray_img[1916]) );
  QDFFS gray_img_reg_15__0__4_ ( .D(n14892), .CK(clk), .Q(gray_img[1924]) );
  QDFFS gray_img_reg_15__1__4_ ( .D(n14891), .CK(clk), .Q(gray_img[1932]) );
  QDFFS gray_img_reg_15__2__4_ ( .D(n14890), .CK(clk), .Q(gray_img[1940]) );
  QDFFS gray_img_reg_15__3__4_ ( .D(n14889), .CK(clk), .Q(gray_img[1948]) );
  QDFFS gray_img_reg_15__4__4_ ( .D(n14888), .CK(clk), .Q(gray_img[1956]) );
  QDFFS gray_img_reg_15__5__4_ ( .D(n14887), .CK(clk), .Q(gray_img[1964]) );
  QDFFS gray_img_reg_15__6__4_ ( .D(n14886), .CK(clk), .Q(gray_img[1972]) );
  QDFFS gray_img_reg_15__7__4_ ( .D(n14885), .CK(clk), .Q(gray_img[1980]) );
  QDFFS gray_img_reg_15__8__4_ ( .D(n14884), .CK(clk), .Q(gray_img[1988]) );
  QDFFS gray_img_reg_15__9__4_ ( .D(n14883), .CK(clk), .Q(gray_img[1996]) );
  QDFFS gray_img_reg_15__10__4_ ( .D(n14882), .CK(clk), .Q(gray_img[2004]) );
  QDFFS gray_img_reg_15__11__4_ ( .D(n14881), .CK(clk), .Q(gray_img[2012]) );
  QDFFS gray_img_reg_15__12__4_ ( .D(n14880), .CK(clk), .Q(gray_img[2020]) );
  QDFFS gray_img_reg_15__13__4_ ( .D(n14879), .CK(clk), .Q(gray_img[2028]) );
  QDFFS gray_img_reg_15__14__4_ ( .D(n14878), .CK(clk), .Q(gray_img[2036]) );
  QDFFS gray_img_reg_15__15__4_ ( .D(n14877), .CK(clk), .Q(gray_img[2044]) );
  QDFFS gray_img_reg_7__1__4_ ( .D(n14871), .CK(clk), .Q(gray_img[908]) );
  QDFFS gray_img_reg_0__4__4_ ( .D(n14253), .CK(clk), .Q(gray_img[36]) );
  QDFFS gray_img_reg_0__5__4_ ( .D(n14244), .CK(clk), .Q(gray_img[44]) );
  QDFFS gray_img_reg_0__6__4_ ( .D(n14235), .CK(clk), .Q(gray_img[52]) );
  QDFFS gray_img_reg_0__7__4_ ( .D(n14226), .CK(clk), .Q(gray_img[60]) );
  QDFFS gray_img_reg_1__4__4_ ( .D(n14209), .CK(clk), .Q(gray_img[164]) );
  QDFFS gray_img_reg_1__5__4_ ( .D(n14200), .CK(clk), .Q(gray_img[172]) );
  QDFFS gray_img_reg_1__6__4_ ( .D(n14191), .CK(clk), .Q(gray_img[180]) );
  QDFFS gray_img_reg_1__7__4_ ( .D(n14182), .CK(clk), .Q(gray_img[188]) );
  QDFFS gray_img_reg_2__4__4_ ( .D(n14165), .CK(clk), .Q(gray_img[292]) );
  QDFFS gray_img_reg_2__5__4_ ( .D(n14156), .CK(clk), .Q(gray_img[300]) );
  QDFFS gray_img_reg_2__6__4_ ( .D(n14147), .CK(clk), .Q(gray_img[308]) );
  QDFFS gray_img_reg_2__7__4_ ( .D(n14138), .CK(clk), .Q(gray_img[316]) );
  QDFFS gray_img_reg_3__4__4_ ( .D(n14121), .CK(clk), .Q(gray_img[420]) );
  QDFFS gray_img_reg_3__5__4_ ( .D(n14112), .CK(clk), .Q(gray_img[428]) );
  QDFFS gray_img_reg_3__6__4_ ( .D(n14103), .CK(clk), .Q(gray_img[436]) );
  QDFFS gray_img_reg_3__7__4_ ( .D(n14094), .CK(clk), .Q(gray_img[444]) );
  QDFFS gray_img_reg_4__0__4_ ( .D(n14069), .CK(clk), .Q(gray_img[516]) );
  QDFFS gray_img_reg_4__1__4_ ( .D(n14060), .CK(clk), .Q(gray_img[524]) );
  QDFFS gray_img_reg_4__2__4_ ( .D(n14051), .CK(clk), .Q(gray_img[532]) );
  QDFFS gray_img_reg_4__3__4_ ( .D(n14042), .CK(clk), .Q(gray_img[540]) );
  QDFFS gray_img_reg_4__4__4_ ( .D(n14033), .CK(clk), .Q(gray_img[548]) );
  QDFFS gray_img_reg_4__5__4_ ( .D(n14024), .CK(clk), .Q(gray_img[556]) );
  QDFFS gray_img_reg_4__6__4_ ( .D(n14015), .CK(clk), .Q(gray_img[564]) );
  QDFFS gray_img_reg_4__7__4_ ( .D(n14006), .CK(clk), .Q(gray_img[572]) );
  QDFFS gray_img_reg_5__0__4_ ( .D(n13981), .CK(clk), .Q(gray_img[644]) );
  QDFFS gray_img_reg_5__1__4_ ( .D(n13972), .CK(clk), .Q(gray_img[652]) );
  QDFFS gray_img_reg_5__2__4_ ( .D(n13963), .CK(clk), .Q(gray_img[660]) );
  QDFFS gray_img_reg_5__3__4_ ( .D(n13955), .CK(clk), .Q(gray_img[668]) );
  QDFFS gray_img_reg_5__4__4_ ( .D(n13947), .CK(clk), .Q(gray_img[676]) );
  QDFFS gray_img_reg_5__5__4_ ( .D(n13940), .CK(clk), .Q(gray_img[684]) );
  QDFFS gray_img_reg_5__6__4_ ( .D(n13933), .CK(clk), .Q(gray_img[692]) );
  QDFFS gray_img_reg_5__7__4_ ( .D(n13927), .CK(clk), .Q(gray_img[700]) );
  QDFFS gray_img_reg_6__0__4_ ( .D(n13905), .CK(clk), .Q(gray_img[772]) );
  QDFFS gray_img_reg_6__1__4_ ( .D(n13899), .CK(clk), .Q(gray_img[780]) );
  QDFFS gray_img_reg_6__2__4_ ( .D(n13893), .CK(clk), .Q(gray_img[788]) );
  QDFFS gray_img_reg_6__3__4_ ( .D(n13887), .CK(clk), .Q(gray_img[796]) );
  QDFFS gray_img_reg_6__4__4_ ( .D(n13881), .CK(clk), .Q(gray_img[804]) );
  QDFFS gray_img_reg_6__5__4_ ( .D(n13875), .CK(clk), .Q(gray_img[812]) );
  QDFFS gray_img_reg_6__6__4_ ( .D(n13869), .CK(clk), .Q(gray_img[820]) );
  QDFFS gray_img_reg_6__7__4_ ( .D(n13863), .CK(clk), .Q(gray_img[828]) );
  QDFFS gray_img_reg_7__0__4_ ( .D(n13841), .CK(clk), .Q(gray_img[900]) );
  QDFFS gray_img_reg_0__2__4_ ( .D(n13798), .CK(clk), .Q(gray_img[20]) );
  QDFFS gray_img_reg_0__3__4_ ( .D(n13788), .CK(clk), .Q(gray_img[28]) );
  QDFFS gray_img_reg_1__2__4_ ( .D(n13768), .CK(clk), .Q(gray_img[148]) );
  QDFFS gray_img_reg_1__3__4_ ( .D(n13758), .CK(clk), .Q(gray_img[156]) );
  QDFFS gray_img_reg_0__1__4_ ( .D(n13750), .CK(clk), .Q(gray_img[12]) );
  QDFFS gray_img_reg_2__0__4_ ( .D(n13732), .CK(clk), .Q(gray_img[260]) );
  QDFFS gray_img_reg_2__1__4_ ( .D(n13703), .CK(clk), .Q(gray_img[268]) );
  QDFFS gray_img_reg_2__2__4_ ( .D(n13677), .CK(clk), .Q(gray_img[276]) );
  QDFFS gray_img_reg_2__3__4_ ( .D(n13654), .CK(clk), .Q(gray_img[284]) );
  QDFFS gray_img_reg_3__0__4_ ( .D(n13634), .CK(clk), .Q(gray_img[388]) );
  QDFFS gray_img_reg_7__2__4_ ( .D(n13630), .CK(clk), .Q(gray_img[916]) );
  QDFFS gray_img_reg_7__3__4_ ( .D(n13629), .CK(clk), .Q(gray_img[924]) );
  QDFFS gray_img_reg_3__1__4_ ( .D(n14874), .CK(clk), .Q(gray_img[396]) );
  QDFFS gray_img_reg_1__0__4_ ( .D(n15069), .CK(clk), .Q(gray_img[132]) );
  QDFFS gray_img_reg_7__4__4_ ( .D(n13628), .CK(clk), .Q(gray_img[932]) );
  QDFFS gray_img_reg_7__5__4_ ( .D(n13627), .CK(clk), .Q(gray_img[940]) );
  QDFFS gray_img_reg_3__2__4_ ( .D(n14873), .CK(clk), .Q(gray_img[404]) );
  QDFFS gray_img_reg_7__6__4_ ( .D(n13626), .CK(clk), .Q(gray_img[948]) );
  QDFFS gray_img_reg_7__7__4_ ( .D(n13625), .CK(clk), .Q(gray_img[956]) );
  QDFFS gray_img_reg_3__3__4_ ( .D(n14872), .CK(clk), .Q(gray_img[412]) );
  QDFFS gray_img_reg_1__1__4_ ( .D(n14875), .CK(clk), .Q(gray_img[140]) );
  QDFFS gray_img_reg_0__0__3_ ( .D(n14677), .CK(clk), .Q(gray_img[3]) );
  QDFFS mem_data_out_reg_shift_0_reg_0__3_ ( .D(n15812), .CK(clk), .Q(
        mem_data_out_reg_shift_0[3]) );
  QDFFS mem_data_out_reg_shift_0_reg_1__3_ ( .D(mem_data_out_reg_shift_0[3]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[11]) );
  QDFFS mem_data_out_reg_shift_0_reg_2__3_ ( .D(mem_data_out_reg_shift_0[11]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[19]) );
  QDFFS mem_data_out_reg_shift_0_reg_3__3_ ( .D(mem_data_out_reg_shift_0[19]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[27]) );
  QDFFS mem_data_out_reg_shift_0_reg_4__3_ ( .D(mem_data_out_reg_shift_0[27]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[35]) );
  QDFFS mem_data_out_reg_shift_0_reg_5__3_ ( .D(mem_data_out_reg_shift_0[35]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[43]) );
  QDFFS mem_data_out_reg_shift_0_reg_6__3_ ( .D(mem_data_out_reg_shift_0[43]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[51]) );
  QDFFS mem_data_out_reg_shift_0_reg_7__3_ ( .D(mem_data_out_reg_shift_0[51]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[59]) );
  QDFFS mem_data_out_reg_shift_0_reg_8__3_ ( .D(mem_data_out_reg_shift_0[59]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[67]) );
  QDFFS mem_data_out_reg_shift_0_reg_9__3_ ( .D(mem_data_out_reg_shift_0[67]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[75]) );
  QDFFS mem_data_out_reg_shift_0_reg_10__3_ ( .D(mem_data_out_reg_shift_0[75]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[83]) );
  QDFFS mem_data_out_reg_shift_0_reg_11__3_ ( .D(mem_data_out_reg_shift_0[83]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[91]) );
  QDFFS mem_data_out_reg_shift_0_reg_12__3_ ( .D(mem_data_out_reg_shift_0[91]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[99]) );
  QDFFS mem_data_out_reg_shift_0_reg_13__3_ ( .D(mem_data_out_reg_shift_0[99]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[107]) );
  QDFFS mem_data_out_reg_shift_0_reg_14__3_ ( .D(mem_data_out_reg_shift_0[107]), .CK(clk), .Q(mem_data_out_reg_shift_0[115]) );
  QDFFS mem_data_out_reg_shift_0_reg_15__3_ ( .D(mem_data_out_reg_shift_0[115]), .CK(clk), .Q(mem_data_out_reg_shift_0[123]) );
  QDFFS mem_data_out_reg_shift_1_reg_0__3_ ( .D(n15829), .CK(clk), .Q(
        mem_data_out_reg_shift_1[3]) );
  QDFFS mem_data_out_reg_shift_1_reg_1__3_ ( .D(mem_data_out_reg_shift_1[3]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[11]) );
  QDFFS mem_data_out_reg_shift_1_reg_3__3_ ( .D(mem_data_out_reg_shift_1[19]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[27]) );
  QDFFS mem_data_out_reg_shift_1_reg_4__3_ ( .D(mem_data_out_reg_shift_1[27]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[35]) );
  QDFFS mem_data_out_reg_shift_1_reg_5__3_ ( .D(mem_data_out_reg_shift_1[35]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[43]) );
  QDFFS mem_data_out_reg_shift_1_reg_6__3_ ( .D(mem_data_out_reg_shift_1[43]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[51]) );
  QDFFS mem_data_out_reg_shift_1_reg_7__3_ ( .D(mem_data_out_reg_shift_1[51]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[59]) );
  QDFFS mem_data_out_reg_shift_1_reg_8__3_ ( .D(mem_data_out_reg_shift_1[59]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[67]) );
  QDFFS mem_data_out_reg_shift_1_reg_9__3_ ( .D(mem_data_out_reg_shift_1[67]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[75]) );
  QDFFS mem_data_out_reg_shift_1_reg_10__3_ ( .D(mem_data_out_reg_shift_1[75]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[83]) );
  QDFFS mem_data_out_reg_shift_1_reg_11__3_ ( .D(mem_data_out_reg_shift_1[83]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[91]) );
  QDFFS mem_data_out_reg_shift_1_reg_12__3_ ( .D(mem_data_out_reg_shift_1[91]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[99]) );
  QDFFS mem_data_out_reg_shift_1_reg_13__3_ ( .D(mem_data_out_reg_shift_1[99]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[107]) );
  QDFFS mem_data_out_reg_shift_1_reg_14__3_ ( .D(mem_data_out_reg_shift_1[107]), .CK(clk), .Q(mem_data_out_reg_shift_1[115]) );
  QDFFS mem_data_out_reg_shift_1_reg_15__3_ ( .D(mem_data_out_reg_shift_1[115]), .CK(clk), .Q(mem_data_out_reg_shift_1[123]) );
  QDFFS mem_data_out_reg_shift_2_reg_0__3_ ( .D(n15837), .CK(clk), .Q(
        mem_data_out_reg_shift_2[3]) );
  QDFFS mem_data_out_reg_shift_2_reg_1__3_ ( .D(mem_data_out_reg_shift_2[3]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[11]) );
  QDFFS mem_data_out_reg_shift_2_reg_2__3_ ( .D(mem_data_out_reg_shift_2[11]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[19]) );
  QDFFS mem_data_out_reg_shift_2_reg_3__3_ ( .D(mem_data_out_reg_shift_2[19]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[27]) );
  QDFFS gray_img_reg_0__8__3_ ( .D(n14869), .CK(clk), .Q(gray_img[67]) );
  QDFFS gray_img_reg_0__9__3_ ( .D(n14868), .CK(clk), .Q(gray_img[75]) );
  QDFFS gray_img_reg_0__10__3_ ( .D(n14867), .CK(clk), .Q(gray_img[83]) );
  QDFFS gray_img_reg_0__11__3_ ( .D(n14866), .CK(clk), .Q(gray_img[91]) );
  QDFFS gray_img_reg_0__12__3_ ( .D(n14865), .CK(clk), .Q(gray_img[99]) );
  QDFFS gray_img_reg_0__13__3_ ( .D(n14864), .CK(clk), .Q(gray_img[107]) );
  QDFFS gray_img_reg_0__14__3_ ( .D(n14863), .CK(clk), .Q(gray_img[115]) );
  QDFFS gray_img_reg_0__15__3_ ( .D(n14862), .CK(clk), .Q(gray_img[123]) );
  QDFFS gray_img_reg_1__8__3_ ( .D(n14861), .CK(clk), .Q(gray_img[195]) );
  QDFFS gray_img_reg_1__9__3_ ( .D(n14860), .CK(clk), .Q(gray_img[203]) );
  QDFFS gray_img_reg_1__10__3_ ( .D(n14859), .CK(clk), .Q(gray_img[211]) );
  QDFFS gray_img_reg_1__11__3_ ( .D(n14858), .CK(clk), .Q(gray_img[219]) );
  QDFFS gray_img_reg_1__12__3_ ( .D(n14857), .CK(clk), .Q(gray_img[227]) );
  QDFFS gray_img_reg_1__13__3_ ( .D(n14856), .CK(clk), .Q(gray_img[235]) );
  QDFFS gray_img_reg_1__14__3_ ( .D(n14855), .CK(clk), .Q(gray_img[243]) );
  QDFFS gray_img_reg_1__15__3_ ( .D(n14854), .CK(clk), .Q(gray_img[251]) );
  QDFFS gray_img_reg_2__8__3_ ( .D(n14853), .CK(clk), .Q(gray_img[323]) );
  QDFFS gray_img_reg_2__9__3_ ( .D(n14852), .CK(clk), .Q(gray_img[331]) );
  QDFFS gray_img_reg_2__10__3_ ( .D(n14851), .CK(clk), .Q(gray_img[339]) );
  QDFFS gray_img_reg_2__11__3_ ( .D(n14850), .CK(clk), .Q(gray_img[347]) );
  QDFFS gray_img_reg_2__12__3_ ( .D(n14849), .CK(clk), .Q(gray_img[355]) );
  QDFFS gray_img_reg_2__13__3_ ( .D(n14848), .CK(clk), .Q(gray_img[363]) );
  QDFFS gray_img_reg_2__14__3_ ( .D(n14847), .CK(clk), .Q(gray_img[371]) );
  QDFFS gray_img_reg_2__15__3_ ( .D(n14846), .CK(clk), .Q(gray_img[379]) );
  QDFFS gray_img_reg_3__8__3_ ( .D(n14845), .CK(clk), .Q(gray_img[451]) );
  QDFFS gray_img_reg_3__9__3_ ( .D(n14844), .CK(clk), .Q(gray_img[459]) );
  QDFFS gray_img_reg_3__10__3_ ( .D(n14843), .CK(clk), .Q(gray_img[467]) );
  QDFFS gray_img_reg_3__11__3_ ( .D(n14842), .CK(clk), .Q(gray_img[475]) );
  QDFFS gray_img_reg_3__12__3_ ( .D(n14841), .CK(clk), .Q(gray_img[483]) );
  QDFFS gray_img_reg_3__13__3_ ( .D(n14840), .CK(clk), .Q(gray_img[491]) );
  QDFFS gray_img_reg_3__14__3_ ( .D(n14839), .CK(clk), .Q(gray_img[499]) );
  QDFFS gray_img_reg_3__15__3_ ( .D(n14838), .CK(clk), .Q(gray_img[507]) );
  QDFFS gray_img_reg_4__8__3_ ( .D(n14837), .CK(clk), .Q(gray_img[579]) );
  QDFFS gray_img_reg_4__9__3_ ( .D(n14836), .CK(clk), .Q(gray_img[587]) );
  QDFFS gray_img_reg_4__10__3_ ( .D(n14835), .CK(clk), .Q(gray_img[595]) );
  QDFFS gray_img_reg_4__11__3_ ( .D(n14834), .CK(clk), .Q(gray_img[603]) );
  QDFFS gray_img_reg_4__12__3_ ( .D(n14833), .CK(clk), .Q(gray_img[611]) );
  QDFFS gray_img_reg_4__13__3_ ( .D(n14832), .CK(clk), .Q(gray_img[619]) );
  QDFFS gray_img_reg_4__14__3_ ( .D(n14831), .CK(clk), .Q(gray_img[627]) );
  QDFFS gray_img_reg_4__15__3_ ( .D(n14830), .CK(clk), .Q(gray_img[635]) );
  QDFFS gray_img_reg_5__8__3_ ( .D(n14829), .CK(clk), .Q(gray_img[707]) );
  QDFFS gray_img_reg_5__9__3_ ( .D(n14828), .CK(clk), .Q(gray_img[715]) );
  QDFFS gray_img_reg_5__10__3_ ( .D(n14827), .CK(clk), .Q(gray_img[723]) );
  QDFFS gray_img_reg_5__11__3_ ( .D(n14826), .CK(clk), .Q(gray_img[731]) );
  QDFFS gray_img_reg_5__12__3_ ( .D(n14825), .CK(clk), .Q(gray_img[739]) );
  QDFFS gray_img_reg_5__13__3_ ( .D(n14824), .CK(clk), .Q(gray_img[747]) );
  QDFFS gray_img_reg_5__14__3_ ( .D(n14823), .CK(clk), .Q(gray_img[755]) );
  QDFFS gray_img_reg_5__15__3_ ( .D(n14822), .CK(clk), .Q(gray_img[763]) );
  QDFFS gray_img_reg_6__8__3_ ( .D(n14821), .CK(clk), .Q(gray_img[835]) );
  QDFFS gray_img_reg_6__9__3_ ( .D(n14820), .CK(clk), .Q(gray_img[843]) );
  QDFFS gray_img_reg_6__10__3_ ( .D(n14819), .CK(clk), .Q(gray_img[851]) );
  QDFFS gray_img_reg_6__11__3_ ( .D(n14818), .CK(clk), .Q(gray_img[859]) );
  QDFFS gray_img_reg_6__12__3_ ( .D(n14817), .CK(clk), .Q(gray_img[867]) );
  QDFFS gray_img_reg_6__13__3_ ( .D(n14816), .CK(clk), .Q(gray_img[875]) );
  QDFFS gray_img_reg_6__14__3_ ( .D(n14815), .CK(clk), .Q(gray_img[883]) );
  QDFFS gray_img_reg_6__15__3_ ( .D(n14814), .CK(clk), .Q(gray_img[891]) );
  QDFFS gray_img_reg_7__8__3_ ( .D(n14813), .CK(clk), .Q(gray_img[963]) );
  QDFFS gray_img_reg_7__9__3_ ( .D(n14812), .CK(clk), .Q(gray_img[971]) );
  QDFFS gray_img_reg_7__10__3_ ( .D(n14811), .CK(clk), .Q(gray_img[979]) );
  QDFFS gray_img_reg_7__11__3_ ( .D(n14810), .CK(clk), .Q(gray_img[987]) );
  QDFFS gray_img_reg_7__12__3_ ( .D(n14809), .CK(clk), .Q(gray_img[995]) );
  QDFFS gray_img_reg_7__13__3_ ( .D(n14808), .CK(clk), .Q(gray_img[1003]) );
  QDFFS gray_img_reg_7__14__3_ ( .D(n14807), .CK(clk), .Q(gray_img[1011]) );
  QDFFS gray_img_reg_7__15__3_ ( .D(n14806), .CK(clk), .Q(gray_img[1019]) );
  QDFFS gray_img_reg_8__0__3_ ( .D(n14805), .CK(clk), .Q(gray_img[1027]) );
  QDFFS gray_img_reg_8__1__3_ ( .D(n14804), .CK(clk), .Q(gray_img[1035]) );
  QDFFS gray_img_reg_8__2__3_ ( .D(n14803), .CK(clk), .Q(gray_img[1043]) );
  QDFFS gray_img_reg_8__3__3_ ( .D(n14802), .CK(clk), .Q(gray_img[1051]) );
  QDFFS gray_img_reg_8__4__3_ ( .D(n14801), .CK(clk), .Q(gray_img[1059]) );
  QDFFS gray_img_reg_8__5__3_ ( .D(n14800), .CK(clk), .Q(gray_img[1067]) );
  QDFFS gray_img_reg_8__6__3_ ( .D(n14799), .CK(clk), .Q(gray_img[1075]) );
  QDFFS gray_img_reg_8__7__3_ ( .D(n14798), .CK(clk), .Q(gray_img[1083]) );
  QDFFS gray_img_reg_8__8__3_ ( .D(n14797), .CK(clk), .Q(gray_img[1091]) );
  QDFFS gray_img_reg_8__9__3_ ( .D(n14796), .CK(clk), .Q(gray_img[1099]) );
  QDFFS gray_img_reg_8__10__3_ ( .D(n14795), .CK(clk), .Q(gray_img[1107]) );
  QDFFS gray_img_reg_8__11__3_ ( .D(n14794), .CK(clk), .Q(gray_img[1115]) );
  QDFFS gray_img_reg_8__12__3_ ( .D(n14793), .CK(clk), .Q(gray_img[1123]) );
  QDFFS gray_img_reg_8__13__3_ ( .D(n14792), .CK(clk), .Q(gray_img[1131]) );
  QDFFS gray_img_reg_8__14__3_ ( .D(n14791), .CK(clk), .Q(gray_img[1139]) );
  QDFFS gray_img_reg_8__15__3_ ( .D(n14790), .CK(clk), .Q(gray_img[1147]) );
  QDFFS gray_img_reg_9__0__3_ ( .D(n14789), .CK(clk), .Q(gray_img[1155]) );
  QDFFS gray_img_reg_9__1__3_ ( .D(n14788), .CK(clk), .Q(gray_img[1163]) );
  QDFFS gray_img_reg_9__2__3_ ( .D(n14787), .CK(clk), .Q(gray_img[1171]) );
  QDFFS gray_img_reg_9__3__3_ ( .D(n14786), .CK(clk), .Q(gray_img[1179]) );
  QDFFS gray_img_reg_9__4__3_ ( .D(n14785), .CK(clk), .Q(gray_img[1187]) );
  QDFFS gray_img_reg_9__5__3_ ( .D(n14784), .CK(clk), .Q(gray_img[1195]) );
  QDFFS gray_img_reg_9__6__3_ ( .D(n14783), .CK(clk), .Q(gray_img[1203]) );
  QDFFS gray_img_reg_9__7__3_ ( .D(n14782), .CK(clk), .Q(gray_img[1211]) );
  QDFFS gray_img_reg_9__8__3_ ( .D(n14781), .CK(clk), .Q(gray_img[1219]) );
  QDFFS gray_img_reg_9__9__3_ ( .D(n14780), .CK(clk), .Q(gray_img[1227]) );
  QDFFS gray_img_reg_9__10__3_ ( .D(n14779), .CK(clk), .Q(gray_img[1235]) );
  QDFFS gray_img_reg_9__11__3_ ( .D(n14778), .CK(clk), .Q(gray_img[1243]) );
  QDFFS gray_img_reg_9__12__3_ ( .D(n14777), .CK(clk), .Q(gray_img[1251]) );
  QDFFS gray_img_reg_9__13__3_ ( .D(n14776), .CK(clk), .Q(gray_img[1259]) );
  QDFFS gray_img_reg_9__14__3_ ( .D(n14775), .CK(clk), .Q(gray_img[1267]) );
  QDFFS gray_img_reg_9__15__3_ ( .D(n14774), .CK(clk), .Q(gray_img[1275]) );
  QDFFS gray_img_reg_10__0__3_ ( .D(n14773), .CK(clk), .Q(gray_img[1283]) );
  QDFFS gray_img_reg_10__1__3_ ( .D(n14772), .CK(clk), .Q(gray_img[1291]) );
  QDFFS gray_img_reg_10__2__3_ ( .D(n14771), .CK(clk), .Q(gray_img[1299]) );
  QDFFS gray_img_reg_10__3__3_ ( .D(n14770), .CK(clk), .Q(gray_img[1307]) );
  QDFFS gray_img_reg_10__4__3_ ( .D(n14769), .CK(clk), .Q(gray_img[1315]) );
  QDFFS gray_img_reg_10__5__3_ ( .D(n14768), .CK(clk), .Q(gray_img[1323]) );
  QDFFS gray_img_reg_10__6__3_ ( .D(n14767), .CK(clk), .Q(gray_img[1331]) );
  QDFFS gray_img_reg_10__7__3_ ( .D(n14766), .CK(clk), .Q(gray_img[1339]) );
  QDFFS gray_img_reg_10__8__3_ ( .D(n14765), .CK(clk), .Q(gray_img[1347]) );
  QDFFS gray_img_reg_10__9__3_ ( .D(n14764), .CK(clk), .Q(gray_img[1355]) );
  QDFFS gray_img_reg_10__10__3_ ( .D(n14763), .CK(clk), .Q(gray_img[1363]) );
  QDFFS gray_img_reg_10__11__3_ ( .D(n14762), .CK(clk), .Q(gray_img[1371]) );
  QDFFS gray_img_reg_10__12__3_ ( .D(n14761), .CK(clk), .Q(gray_img[1379]) );
  QDFFS gray_img_reg_10__13__3_ ( .D(n14760), .CK(clk), .Q(gray_img[1387]) );
  QDFFS gray_img_reg_10__14__3_ ( .D(n14759), .CK(clk), .Q(gray_img[1395]) );
  QDFFS gray_img_reg_10__15__3_ ( .D(n14758), .CK(clk), .Q(gray_img[1403]) );
  QDFFS gray_img_reg_11__0__3_ ( .D(n14757), .CK(clk), .Q(gray_img[1411]) );
  QDFFS gray_img_reg_11__1__3_ ( .D(n14756), .CK(clk), .Q(gray_img[1419]) );
  QDFFS gray_img_reg_11__2__3_ ( .D(n14755), .CK(clk), .Q(gray_img[1427]) );
  QDFFS gray_img_reg_11__3__3_ ( .D(n14754), .CK(clk), .Q(gray_img[1435]) );
  QDFFS gray_img_reg_11__4__3_ ( .D(n14753), .CK(clk), .Q(gray_img[1443]) );
  QDFFS gray_img_reg_11__5__3_ ( .D(n14752), .CK(clk), .Q(gray_img[1451]) );
  QDFFS gray_img_reg_11__6__3_ ( .D(n14751), .CK(clk), .Q(gray_img[1459]) );
  QDFFS gray_img_reg_11__7__3_ ( .D(n14750), .CK(clk), .Q(gray_img[1467]) );
  QDFFS gray_img_reg_11__8__3_ ( .D(n14749), .CK(clk), .Q(gray_img[1475]) );
  QDFFS gray_img_reg_11__9__3_ ( .D(n14748), .CK(clk), .Q(gray_img[1483]) );
  QDFFS gray_img_reg_11__10__3_ ( .D(n14747), .CK(clk), .Q(gray_img[1491]) );
  QDFFS gray_img_reg_11__11__3_ ( .D(n14746), .CK(clk), .Q(gray_img[1499]) );
  QDFFS gray_img_reg_11__12__3_ ( .D(n14745), .CK(clk), .Q(gray_img[1507]) );
  QDFFS gray_img_reg_11__13__3_ ( .D(n14744), .CK(clk), .Q(gray_img[1515]) );
  QDFFS gray_img_reg_11__14__3_ ( .D(n14743), .CK(clk), .Q(gray_img[1523]) );
  QDFFS gray_img_reg_11__15__3_ ( .D(n14742), .CK(clk), .Q(gray_img[1531]) );
  QDFFS gray_img_reg_12__0__3_ ( .D(n14741), .CK(clk), .Q(gray_img[1539]) );
  QDFFS gray_img_reg_12__1__3_ ( .D(n14740), .CK(clk), .Q(gray_img[1547]) );
  QDFFS gray_img_reg_12__2__3_ ( .D(n14739), .CK(clk), .Q(gray_img[1555]) );
  QDFFS gray_img_reg_12__3__3_ ( .D(n14738), .CK(clk), .Q(gray_img[1563]) );
  QDFFS gray_img_reg_12__4__3_ ( .D(n14737), .CK(clk), .Q(gray_img[1571]) );
  QDFFS gray_img_reg_12__5__3_ ( .D(n14736), .CK(clk), .Q(gray_img[1579]) );
  QDFFS gray_img_reg_12__6__3_ ( .D(n14735), .CK(clk), .Q(gray_img[1587]) );
  QDFFS gray_img_reg_12__7__3_ ( .D(n14734), .CK(clk), .Q(gray_img[1595]) );
  QDFFS gray_img_reg_12__8__3_ ( .D(n14733), .CK(clk), .Q(gray_img[1603]) );
  QDFFS gray_img_reg_12__9__3_ ( .D(n14732), .CK(clk), .Q(gray_img[1611]) );
  QDFFS gray_img_reg_12__10__3_ ( .D(n14731), .CK(clk), .Q(gray_img[1619]) );
  QDFFS gray_img_reg_12__11__3_ ( .D(n14730), .CK(clk), .Q(gray_img[1627]) );
  QDFFS gray_img_reg_12__12__3_ ( .D(n14729), .CK(clk), .Q(gray_img[1635]) );
  QDFFS gray_img_reg_12__13__3_ ( .D(n14728), .CK(clk), .Q(gray_img[1643]) );
  QDFFS gray_img_reg_12__14__3_ ( .D(n14727), .CK(clk), .Q(gray_img[1651]) );
  QDFFS gray_img_reg_12__15__3_ ( .D(n14726), .CK(clk), .Q(gray_img[1659]) );
  QDFFS gray_img_reg_13__0__3_ ( .D(n14725), .CK(clk), .Q(gray_img[1667]) );
  QDFFS gray_img_reg_13__1__3_ ( .D(n14724), .CK(clk), .Q(gray_img[1675]) );
  QDFFS gray_img_reg_13__2__3_ ( .D(n14723), .CK(clk), .Q(gray_img[1683]) );
  QDFFS gray_img_reg_13__3__3_ ( .D(n14722), .CK(clk), .Q(gray_img[1691]) );
  QDFFS gray_img_reg_13__4__3_ ( .D(n14721), .CK(clk), .Q(gray_img[1699]) );
  QDFFS gray_img_reg_13__5__3_ ( .D(n14720), .CK(clk), .Q(gray_img[1707]) );
  QDFFS gray_img_reg_13__6__3_ ( .D(n14719), .CK(clk), .Q(gray_img[1715]) );
  QDFFS gray_img_reg_13__7__3_ ( .D(n14718), .CK(clk), .Q(gray_img[1723]) );
  QDFFS gray_img_reg_13__8__3_ ( .D(n14717), .CK(clk), .Q(gray_img[1731]) );
  QDFFS gray_img_reg_13__9__3_ ( .D(n14716), .CK(clk), .Q(gray_img[1739]) );
  QDFFS gray_img_reg_13__10__3_ ( .D(n14715), .CK(clk), .Q(gray_img[1747]) );
  QDFFS gray_img_reg_13__11__3_ ( .D(n14714), .CK(clk), .Q(gray_img[1755]) );
  QDFFS gray_img_reg_13__12__3_ ( .D(n14713), .CK(clk), .Q(gray_img[1763]) );
  QDFFS gray_img_reg_13__13__3_ ( .D(n14712), .CK(clk), .Q(gray_img[1771]) );
  QDFFS gray_img_reg_13__14__3_ ( .D(n14711), .CK(clk), .Q(gray_img[1779]) );
  QDFFS gray_img_reg_13__15__3_ ( .D(n14710), .CK(clk), .Q(gray_img[1787]) );
  QDFFS gray_img_reg_14__0__3_ ( .D(n14709), .CK(clk), .Q(gray_img[1795]) );
  QDFFS gray_img_reg_14__1__3_ ( .D(n14708), .CK(clk), .Q(gray_img[1803]) );
  QDFFS gray_img_reg_14__2__3_ ( .D(n14707), .CK(clk), .Q(gray_img[1811]) );
  QDFFS gray_img_reg_14__3__3_ ( .D(n14706), .CK(clk), .Q(gray_img[1819]) );
  QDFFS gray_img_reg_14__4__3_ ( .D(n14705), .CK(clk), .Q(gray_img[1827]) );
  QDFFS gray_img_reg_14__5__3_ ( .D(n14704), .CK(clk), .Q(gray_img[1835]) );
  QDFFS gray_img_reg_14__6__3_ ( .D(n14703), .CK(clk), .Q(gray_img[1843]) );
  QDFFS gray_img_reg_14__7__3_ ( .D(n14702), .CK(clk), .Q(gray_img[1851]) );
  QDFFS gray_img_reg_14__8__3_ ( .D(n14701), .CK(clk), .Q(gray_img[1859]) );
  QDFFS gray_img_reg_14__9__3_ ( .D(n14700), .CK(clk), .Q(gray_img[1867]) );
  QDFFS gray_img_reg_14__10__3_ ( .D(n14699), .CK(clk), .Q(gray_img[1875]) );
  QDFFS gray_img_reg_14__11__3_ ( .D(n14698), .CK(clk), .Q(gray_img[1883]) );
  QDFFS gray_img_reg_14__12__3_ ( .D(n14697), .CK(clk), .Q(gray_img[1891]) );
  QDFFS gray_img_reg_14__13__3_ ( .D(n14696), .CK(clk), .Q(gray_img[1899]) );
  QDFFS gray_img_reg_14__14__3_ ( .D(n14695), .CK(clk), .Q(gray_img[1907]) );
  QDFFS gray_img_reg_14__15__3_ ( .D(n14694), .CK(clk), .Q(gray_img[1915]) );
  QDFFS gray_img_reg_15__0__3_ ( .D(n14693), .CK(clk), .Q(gray_img[1923]) );
  QDFFS gray_img_reg_15__1__3_ ( .D(n14692), .CK(clk), .Q(gray_img[1931]) );
  QDFFS gray_img_reg_15__2__3_ ( .D(n14691), .CK(clk), .Q(gray_img[1939]) );
  QDFFS gray_img_reg_15__3__3_ ( .D(n14690), .CK(clk), .Q(gray_img[1947]) );
  QDFFS gray_img_reg_15__4__3_ ( .D(n14689), .CK(clk), .Q(gray_img[1955]) );
  QDFFS gray_img_reg_15__5__3_ ( .D(n14688), .CK(clk), .Q(gray_img[1963]) );
  QDFFS gray_img_reg_15__6__3_ ( .D(n14687), .CK(clk), .Q(gray_img[1971]) );
  QDFFS gray_img_reg_15__7__3_ ( .D(n14686), .CK(clk), .Q(gray_img[1979]) );
  QDFFS gray_img_reg_15__8__3_ ( .D(n14685), .CK(clk), .Q(gray_img[1987]) );
  QDFFS gray_img_reg_15__9__3_ ( .D(n14684), .CK(clk), .Q(gray_img[1995]) );
  QDFFS gray_img_reg_15__10__3_ ( .D(n14683), .CK(clk), .Q(gray_img[2003]) );
  QDFFS gray_img_reg_15__11__3_ ( .D(n14682), .CK(clk), .Q(gray_img[2011]) );
  QDFFS gray_img_reg_15__12__3_ ( .D(n14681), .CK(clk), .Q(gray_img[2019]) );
  QDFFS gray_img_reg_15__13__3_ ( .D(n14680), .CK(clk), .Q(gray_img[2027]) );
  QDFFS gray_img_reg_15__14__3_ ( .D(n14679), .CK(clk), .Q(gray_img[2035]) );
  QDFFS gray_img_reg_15__15__3_ ( .D(n14678), .CK(clk), .Q(gray_img[2043]) );
  QDFFS gray_img_reg_5__7__3_ ( .D(n14671), .CK(clk), .Q(gray_img[699]) );
  QDFFS gray_img_reg_0__4__3_ ( .D(n14254), .CK(clk), .Q(gray_img[35]) );
  QDFFS gray_img_reg_0__5__3_ ( .D(n14245), .CK(clk), .Q(gray_img[43]) );
  QDFFS gray_img_reg_0__6__3_ ( .D(n14236), .CK(clk), .Q(gray_img[51]) );
  QDFFS gray_img_reg_0__7__3_ ( .D(n14227), .CK(clk), .Q(gray_img[59]) );
  QDFFS gray_img_reg_1__4__3_ ( .D(n14210), .CK(clk), .Q(gray_img[163]) );
  QDFFS gray_img_reg_1__5__3_ ( .D(n14201), .CK(clk), .Q(gray_img[171]) );
  QDFFS gray_img_reg_1__6__3_ ( .D(n14192), .CK(clk), .Q(gray_img[179]) );
  QDFFS gray_img_reg_1__7__3_ ( .D(n14183), .CK(clk), .Q(gray_img[187]) );
  QDFFS gray_img_reg_2__4__3_ ( .D(n14166), .CK(clk), .Q(gray_img[291]) );
  QDFFS gray_img_reg_2__5__3_ ( .D(n14157), .CK(clk), .Q(gray_img[299]) );
  QDFFS gray_img_reg_2__6__3_ ( .D(n14148), .CK(clk), .Q(gray_img[307]) );
  QDFFS gray_img_reg_2__7__3_ ( .D(n14139), .CK(clk), .Q(gray_img[315]) );
  QDFFS gray_img_reg_3__4__3_ ( .D(n14122), .CK(clk), .Q(gray_img[419]) );
  QDFFS gray_img_reg_3__5__3_ ( .D(n14113), .CK(clk), .Q(gray_img[427]) );
  QDFFS gray_img_reg_3__6__3_ ( .D(n14104), .CK(clk), .Q(gray_img[435]) );
  QDFFS gray_img_reg_3__7__3_ ( .D(n14095), .CK(clk), .Q(gray_img[443]) );
  QDFFS gray_img_reg_4__0__3_ ( .D(n14070), .CK(clk), .Q(gray_img[515]) );
  QDFFS gray_img_reg_4__1__3_ ( .D(n14061), .CK(clk), .Q(gray_img[523]) );
  QDFFS gray_img_reg_4__2__3_ ( .D(n14052), .CK(clk), .Q(gray_img[531]) );
  QDFFS gray_img_reg_4__3__3_ ( .D(n14043), .CK(clk), .Q(gray_img[539]) );
  QDFFS gray_img_reg_4__4__3_ ( .D(n14034), .CK(clk), .Q(gray_img[547]) );
  QDFFS gray_img_reg_4__5__3_ ( .D(n14025), .CK(clk), .Q(gray_img[555]) );
  QDFFS gray_img_reg_4__6__3_ ( .D(n14016), .CK(clk), .Q(gray_img[563]) );
  QDFFS gray_img_reg_4__7__3_ ( .D(n14007), .CK(clk), .Q(gray_img[571]) );
  QDFFS gray_img_reg_5__0__3_ ( .D(n13982), .CK(clk), .Q(gray_img[643]) );
  QDFFS gray_img_reg_5__1__3_ ( .D(n13973), .CK(clk), .Q(gray_img[651]) );
  QDFFS gray_img_reg_5__2__3_ ( .D(n13964), .CK(clk), .Q(gray_img[659]) );
  QDFFS gray_img_reg_5__3__3_ ( .D(n13956), .CK(clk), .Q(gray_img[667]) );
  QDFFS gray_img_reg_5__4__3_ ( .D(n13948), .CK(clk), .Q(gray_img[675]) );
  QDFFS gray_img_reg_5__5__3_ ( .D(n13941), .CK(clk), .Q(gray_img[683]) );
  QDFFS gray_img_reg_5__6__3_ ( .D(n13934), .CK(clk), .Q(gray_img[691]) );
  QDFFS gray_img_reg_0__2__3_ ( .D(n13799), .CK(clk), .Q(gray_img[19]) );
  QDFFS gray_img_reg_0__3__3_ ( .D(n13789), .CK(clk), .Q(gray_img[27]) );
  QDFFS gray_img_reg_1__2__3_ ( .D(n13769), .CK(clk), .Q(gray_img[147]) );
  QDFFS gray_img_reg_1__3__3_ ( .D(n13759), .CK(clk), .Q(gray_img[155]) );
  QDFFS gray_img_reg_0__1__3_ ( .D(n13751), .CK(clk), .Q(gray_img[11]) );
  QDFFS gray_img_reg_2__0__3_ ( .D(n13733), .CK(clk), .Q(gray_img[259]) );
  QDFFS gray_img_reg_2__1__3_ ( .D(n13704), .CK(clk), .Q(gray_img[267]) );
  QDFFS gray_img_reg_2__2__3_ ( .D(n13678), .CK(clk), .Q(gray_img[275]) );
  QDFFS gray_img_reg_2__3__3_ ( .D(n13655), .CK(clk), .Q(gray_img[283]) );
  QDFFS gray_img_reg_6__0__3_ ( .D(n13650), .CK(clk), .Q(gray_img[771]) );
  QDFFS gray_img_reg_6__1__3_ ( .D(n13649), .CK(clk), .Q(gray_img[779]) );
  QDFFS gray_img_reg_6__2__3_ ( .D(n13648), .CK(clk), .Q(gray_img[787]) );
  QDFFS gray_img_reg_6__3__3_ ( .D(n13647), .CK(clk), .Q(gray_img[795]) );
  QDFFS gray_img_reg_6__4__3_ ( .D(n13646), .CK(clk), .Q(gray_img[803]) );
  QDFFS gray_img_reg_6__5__3_ ( .D(n13645), .CK(clk), .Q(gray_img[811]) );
  QDFFS gray_img_reg_6__6__3_ ( .D(n13644), .CK(clk), .Q(gray_img[819]) );
  QDFFS gray_img_reg_6__7__3_ ( .D(n13643), .CK(clk), .Q(gray_img[827]) );
  QDFFS gray_img_reg_7__0__3_ ( .D(n13642), .CK(clk), .Q(gray_img[899]) );
  QDFFS gray_img_reg_7__1__3_ ( .D(n13641), .CK(clk), .Q(gray_img[907]) );
  QDFFS gray_img_reg_3__0__3_ ( .D(n14870), .CK(clk), .Q(gray_img[387]) );
  QDFFS gray_img_reg_7__2__3_ ( .D(n13640), .CK(clk), .Q(gray_img[915]) );
  QDFFS gray_img_reg_7__3__3_ ( .D(n13639), .CK(clk), .Q(gray_img[923]) );
  QDFFS gray_img_reg_3__1__3_ ( .D(n14674), .CK(clk), .Q(gray_img[395]) );
  QDFFS gray_img_reg_1__0__3_ ( .D(n14676), .CK(clk), .Q(gray_img[131]) );
  QDFFS gray_img_reg_7__4__3_ ( .D(n13638), .CK(clk), .Q(gray_img[931]) );
  QDFFS gray_img_reg_7__5__3_ ( .D(n13637), .CK(clk), .Q(gray_img[939]) );
  QDFFS gray_img_reg_3__2__3_ ( .D(n14673), .CK(clk), .Q(gray_img[403]) );
  QDFFS gray_img_reg_7__6__3_ ( .D(n13636), .CK(clk), .Q(gray_img[947]) );
  QDFFS gray_img_reg_7__7__3_ ( .D(n13635), .CK(clk), .Q(gray_img[955]) );
  QDFFS gray_img_reg_3__3__3_ ( .D(n14672), .CK(clk), .Q(gray_img[411]) );
  QDFFS gray_img_reg_1__1__3_ ( .D(n14675), .CK(clk), .Q(gray_img[139]) );
  QDFFS gray_img_reg_0__0__2_ ( .D(n14477), .CK(clk), .Q(gray_img[2]) );
  QDFFS mem_data_out_reg_shift_0_reg_0__2_ ( .D(n15813), .CK(clk), .Q(
        mem_data_out_reg_shift_0[2]) );
  QDFFS mem_data_out_reg_shift_0_reg_1__2_ ( .D(mem_data_out_reg_shift_0[2]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[10]) );
  QDFFS mem_data_out_reg_shift_0_reg_2__2_ ( .D(mem_data_out_reg_shift_0[10]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[18]) );
  QDFFS mem_data_out_reg_shift_0_reg_3__2_ ( .D(mem_data_out_reg_shift_0[18]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[26]) );
  QDFFS mem_data_out_reg_shift_0_reg_4__2_ ( .D(mem_data_out_reg_shift_0[26]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[34]) );
  QDFFS mem_data_out_reg_shift_0_reg_5__2_ ( .D(mem_data_out_reg_shift_0[34]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[42]) );
  QDFFS mem_data_out_reg_shift_0_reg_6__2_ ( .D(mem_data_out_reg_shift_0[42]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[50]) );
  QDFFS mem_data_out_reg_shift_0_reg_7__2_ ( .D(mem_data_out_reg_shift_0[50]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[58]) );
  QDFFS mem_data_out_reg_shift_0_reg_8__2_ ( .D(mem_data_out_reg_shift_0[58]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[66]) );
  QDFFS mem_data_out_reg_shift_0_reg_9__2_ ( .D(mem_data_out_reg_shift_0[66]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[74]) );
  QDFFS mem_data_out_reg_shift_0_reg_10__2_ ( .D(mem_data_out_reg_shift_0[74]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[82]) );
  QDFFS mem_data_out_reg_shift_0_reg_11__2_ ( .D(mem_data_out_reg_shift_0[82]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[90]) );
  QDFFS mem_data_out_reg_shift_0_reg_12__2_ ( .D(mem_data_out_reg_shift_0[90]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[98]) );
  QDFFS mem_data_out_reg_shift_0_reg_13__2_ ( .D(mem_data_out_reg_shift_0[98]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[106]) );
  QDFFS mem_data_out_reg_shift_0_reg_14__2_ ( .D(mem_data_out_reg_shift_0[106]), .CK(clk), .Q(mem_data_out_reg_shift_0[114]) );
  QDFFS mem_data_out_reg_shift_0_reg_15__2_ ( .D(mem_data_out_reg_shift_0[114]), .CK(clk), .Q(mem_data_out_reg_shift_0[122]) );
  QDFFS mem_data_out_reg_shift_1_reg_0__2_ ( .D(n15830), .CK(clk), .Q(
        mem_data_out_reg_shift_1[2]) );
  QDFFS mem_data_out_reg_shift_1_reg_1__2_ ( .D(mem_data_out_reg_shift_1[2]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[10]) );
  QDFFS mem_data_out_reg_shift_1_reg_3__2_ ( .D(mem_data_out_reg_shift_1[18]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[26]) );
  QDFFS mem_data_out_reg_shift_1_reg_4__2_ ( .D(mem_data_out_reg_shift_1[26]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[34]) );
  QDFFS mem_data_out_reg_shift_1_reg_5__2_ ( .D(mem_data_out_reg_shift_1[34]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[42]) );
  QDFFS mem_data_out_reg_shift_1_reg_6__2_ ( .D(mem_data_out_reg_shift_1[42]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[50]) );
  QDFFS mem_data_out_reg_shift_1_reg_7__2_ ( .D(mem_data_out_reg_shift_1[50]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[58]) );
  QDFFS mem_data_out_reg_shift_1_reg_8__2_ ( .D(mem_data_out_reg_shift_1[58]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[66]) );
  QDFFS mem_data_out_reg_shift_1_reg_9__2_ ( .D(mem_data_out_reg_shift_1[66]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[74]) );
  QDFFS mem_data_out_reg_shift_1_reg_10__2_ ( .D(mem_data_out_reg_shift_1[74]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[82]) );
  QDFFS mem_data_out_reg_shift_1_reg_11__2_ ( .D(mem_data_out_reg_shift_1[82]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[90]) );
  QDFFS mem_data_out_reg_shift_1_reg_12__2_ ( .D(mem_data_out_reg_shift_1[90]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[98]) );
  QDFFS mem_data_out_reg_shift_1_reg_13__2_ ( .D(mem_data_out_reg_shift_1[98]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[106]) );
  QDFFS mem_data_out_reg_shift_1_reg_14__2_ ( .D(mem_data_out_reg_shift_1[106]), .CK(clk), .Q(mem_data_out_reg_shift_1[114]) );
  QDFFS mem_data_out_reg_shift_1_reg_15__2_ ( .D(mem_data_out_reg_shift_1[114]), .CK(clk), .Q(mem_data_out_reg_shift_1[122]) );
  QDFFS mem_data_out_reg_shift_2_reg_0__2_ ( .D(n15838), .CK(clk), .Q(
        mem_data_out_reg_shift_2[2]) );
  QDFFS mem_data_out_reg_shift_2_reg_1__2_ ( .D(mem_data_out_reg_shift_2[2]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[10]) );
  QDFFS mem_data_out_reg_shift_2_reg_2__2_ ( .D(mem_data_out_reg_shift_2[10]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[18]) );
  QDFFS mem_data_out_reg_shift_2_reg_3__2_ ( .D(mem_data_out_reg_shift_2[18]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[26]) );
  QDFFS gray_img_reg_0__8__2_ ( .D(n14669), .CK(clk), .Q(gray_img[66]) );
  QDFFS gray_img_reg_0__9__2_ ( .D(n14668), .CK(clk), .Q(gray_img[74]) );
  QDFFS gray_img_reg_0__10__2_ ( .D(n14667), .CK(clk), .Q(gray_img[82]) );
  QDFFS gray_img_reg_0__11__2_ ( .D(n14666), .CK(clk), .Q(gray_img[90]) );
  QDFFS gray_img_reg_0__12__2_ ( .D(n14665), .CK(clk), .Q(gray_img[98]) );
  QDFFS gray_img_reg_0__13__2_ ( .D(n14664), .CK(clk), .Q(gray_img[106]) );
  QDFFS gray_img_reg_0__14__2_ ( .D(n14663), .CK(clk), .Q(gray_img[114]) );
  QDFFS gray_img_reg_0__15__2_ ( .D(n14662), .CK(clk), .Q(gray_img[122]) );
  QDFFS gray_img_reg_1__8__2_ ( .D(n14661), .CK(clk), .Q(gray_img[194]) );
  QDFFS gray_img_reg_1__9__2_ ( .D(n14660), .CK(clk), .Q(gray_img[202]) );
  QDFFS gray_img_reg_1__10__2_ ( .D(n14659), .CK(clk), .Q(gray_img[210]) );
  QDFFS gray_img_reg_1__11__2_ ( .D(n14658), .CK(clk), .Q(gray_img[218]) );
  QDFFS gray_img_reg_1__12__2_ ( .D(n14657), .CK(clk), .Q(gray_img[226]) );
  QDFFS gray_img_reg_1__13__2_ ( .D(n14656), .CK(clk), .Q(gray_img[234]) );
  QDFFS gray_img_reg_1__14__2_ ( .D(n14655), .CK(clk), .Q(gray_img[242]) );
  QDFFS gray_img_reg_1__15__2_ ( .D(n14654), .CK(clk), .Q(gray_img[250]) );
  QDFFS gray_img_reg_2__8__2_ ( .D(n14653), .CK(clk), .Q(gray_img[322]) );
  QDFFS gray_img_reg_2__9__2_ ( .D(n14652), .CK(clk), .Q(gray_img[330]) );
  QDFFS gray_img_reg_2__10__2_ ( .D(n14651), .CK(clk), .Q(gray_img[338]) );
  QDFFS gray_img_reg_2__11__2_ ( .D(n14650), .CK(clk), .Q(gray_img[346]) );
  QDFFS gray_img_reg_2__12__2_ ( .D(n14649), .CK(clk), .Q(gray_img[354]) );
  QDFFS gray_img_reg_2__13__2_ ( .D(n14648), .CK(clk), .Q(gray_img[362]) );
  QDFFS gray_img_reg_2__14__2_ ( .D(n14647), .CK(clk), .Q(gray_img[370]) );
  QDFFS gray_img_reg_2__15__2_ ( .D(n14646), .CK(clk), .Q(gray_img[378]) );
  QDFFS gray_img_reg_3__9__2_ ( .D(n14644), .CK(clk), .Q(gray_img[458]) );
  QDFFS gray_img_reg_3__10__2_ ( .D(n14643), .CK(clk), .Q(gray_img[466]) );
  QDFFS gray_img_reg_3__11__2_ ( .D(n14642), .CK(clk), .Q(gray_img[474]) );
  QDFFS gray_img_reg_3__12__2_ ( .D(n14641), .CK(clk), .Q(gray_img[482]) );
  QDFFS gray_img_reg_3__13__2_ ( .D(n14640), .CK(clk), .Q(gray_img[490]) );
  QDFFS gray_img_reg_3__14__2_ ( .D(n14639), .CK(clk), .Q(gray_img[498]) );
  QDFFS gray_img_reg_3__15__2_ ( .D(n14638), .CK(clk), .Q(gray_img[506]) );
  QDFFS gray_img_reg_4__8__2_ ( .D(n14637), .CK(clk), .Q(gray_img[578]) );
  QDFFS gray_img_reg_4__9__2_ ( .D(n14636), .CK(clk), .Q(gray_img[586]) );
  QDFFS gray_img_reg_4__10__2_ ( .D(n14635), .CK(clk), .Q(gray_img[594]) );
  QDFFS gray_img_reg_4__11__2_ ( .D(n14634), .CK(clk), .Q(gray_img[602]) );
  QDFFS gray_img_reg_4__12__2_ ( .D(n14633), .CK(clk), .Q(gray_img[610]) );
  QDFFS gray_img_reg_4__13__2_ ( .D(n14632), .CK(clk), .Q(gray_img[618]) );
  QDFFS gray_img_reg_4__14__2_ ( .D(n14631), .CK(clk), .Q(gray_img[626]) );
  QDFFS gray_img_reg_4__15__2_ ( .D(n14630), .CK(clk), .Q(gray_img[634]) );
  QDFFS gray_img_reg_5__8__2_ ( .D(n14629), .CK(clk), .Q(gray_img[706]) );
  QDFFS gray_img_reg_5__9__2_ ( .D(n14628), .CK(clk), .Q(gray_img[714]) );
  QDFFS gray_img_reg_5__10__2_ ( .D(n14627), .CK(clk), .Q(gray_img[722]) );
  QDFFS gray_img_reg_5__11__2_ ( .D(n14626), .CK(clk), .Q(gray_img[730]) );
  QDFFS gray_img_reg_5__12__2_ ( .D(n14625), .CK(clk), .Q(gray_img[738]) );
  QDFFS gray_img_reg_5__13__2_ ( .D(n14624), .CK(clk), .Q(gray_img[746]) );
  QDFFS gray_img_reg_5__14__2_ ( .D(n14623), .CK(clk), .Q(gray_img[754]) );
  QDFFS gray_img_reg_5__15__2_ ( .D(n14622), .CK(clk), .Q(gray_img[762]) );
  QDFFS gray_img_reg_6__8__2_ ( .D(n14621), .CK(clk), .Q(gray_img[834]) );
  QDFFS gray_img_reg_6__9__2_ ( .D(n14620), .CK(clk), .Q(gray_img[842]) );
  QDFFS gray_img_reg_6__12__2_ ( .D(n14617), .CK(clk), .Q(gray_img[866]) );
  QDFFS gray_img_reg_6__13__2_ ( .D(n14616), .CK(clk), .Q(gray_img[874]) );
  QDFFS gray_img_reg_6__14__2_ ( .D(n14615), .CK(clk), .Q(gray_img[882]) );
  QDFFS gray_img_reg_6__15__2_ ( .D(n14614), .CK(clk), .Q(gray_img[890]) );
  QDFFS gray_img_reg_7__8__2_ ( .D(n14613), .CK(clk), .Q(gray_img[962]) );
  QDFFS gray_img_reg_7__9__2_ ( .D(n14612), .CK(clk), .Q(gray_img[970]) );
  QDFFS gray_img_reg_7__10__2_ ( .D(n14611), .CK(clk), .Q(gray_img[978]) );
  QDFFS gray_img_reg_7__11__2_ ( .D(n14610), .CK(clk), .Q(gray_img[986]) );
  QDFFS gray_img_reg_7__12__2_ ( .D(n14609), .CK(clk), .Q(gray_img[994]) );
  QDFFS gray_img_reg_7__13__2_ ( .D(n14608), .CK(clk), .Q(gray_img[1002]) );
  QDFFS gray_img_reg_7__14__2_ ( .D(n14607), .CK(clk), .Q(gray_img[1010]) );
  QDFFS gray_img_reg_7__15__2_ ( .D(n14606), .CK(clk), .Q(gray_img[1018]) );
  QDFFS gray_img_reg_8__0__2_ ( .D(n14605), .CK(clk), .Q(gray_img[1026]) );
  QDFFS gray_img_reg_8__2__2_ ( .D(n14603), .CK(clk), .Q(gray_img[1042]) );
  QDFFS gray_img_reg_8__3__2_ ( .D(n14602), .CK(clk), .Q(gray_img[1050]) );
  QDFFS gray_img_reg_8__4__2_ ( .D(n14601), .CK(clk), .Q(gray_img[1058]) );
  QDFFS gray_img_reg_8__5__2_ ( .D(n14600), .CK(clk), .Q(gray_img[1066]) );
  QDFFS gray_img_reg_8__6__2_ ( .D(n14599), .CK(clk), .Q(gray_img[1074]) );
  QDFFS gray_img_reg_8__7__2_ ( .D(n14598), .CK(clk), .Q(gray_img[1082]) );
  QDFFS gray_img_reg_8__8__2_ ( .D(n14597), .CK(clk), .Q(gray_img[1090]) );
  QDFFS gray_img_reg_8__9__2_ ( .D(n14596), .CK(clk), .Q(gray_img[1098]) );
  QDFFS gray_img_reg_8__10__2_ ( .D(n14595), .CK(clk), .Q(gray_img[1106]) );
  QDFFS gray_img_reg_8__11__2_ ( .D(n14594), .CK(clk), .Q(gray_img[1114]) );
  QDFFS gray_img_reg_8__12__2_ ( .D(n14593), .CK(clk), .Q(gray_img[1122]) );
  QDFFS gray_img_reg_8__13__2_ ( .D(n14592), .CK(clk), .Q(gray_img[1130]) );
  QDFFS gray_img_reg_8__14__2_ ( .D(n14591), .CK(clk), .Q(gray_img[1138]) );
  QDFFS gray_img_reg_8__15__2_ ( .D(n14590), .CK(clk), .Q(gray_img[1146]) );
  QDFFS gray_img_reg_9__0__2_ ( .D(n14589), .CK(clk), .Q(gray_img[1154]) );
  QDFFS gray_img_reg_9__1__2_ ( .D(n14588), .CK(clk), .Q(gray_img[1162]) );
  QDFFS gray_img_reg_9__4__2_ ( .D(n14585), .CK(clk), .Q(gray_img[1186]) );
  QDFFS gray_img_reg_9__5__2_ ( .D(n14584), .CK(clk), .Q(gray_img[1194]) );
  QDFFS gray_img_reg_9__6__2_ ( .D(n14583), .CK(clk), .Q(gray_img[1202]) );
  QDFFS gray_img_reg_9__7__2_ ( .D(n14582), .CK(clk), .Q(gray_img[1210]) );
  QDFFS gray_img_reg_9__8__2_ ( .D(n14581), .CK(clk), .Q(gray_img[1218]) );
  QDFFS gray_img_reg_9__9__2_ ( .D(n14580), .CK(clk), .Q(gray_img[1226]) );
  QDFFS gray_img_reg_9__10__2_ ( .D(n14579), .CK(clk), .Q(gray_img[1234]) );
  QDFFS gray_img_reg_9__11__2_ ( .D(n14578), .CK(clk), .Q(gray_img[1242]) );
  QDFFS gray_img_reg_9__12__2_ ( .D(n14577), .CK(clk), .Q(gray_img[1250]) );
  QDFFS gray_img_reg_9__13__2_ ( .D(n14576), .CK(clk), .Q(gray_img[1258]) );
  QDFFS gray_img_reg_9__14__2_ ( .D(n14575), .CK(clk), .Q(gray_img[1266]) );
  QDFFS gray_img_reg_9__15__2_ ( .D(n14574), .CK(clk), .Q(gray_img[1274]) );
  QDFFS gray_img_reg_10__0__2_ ( .D(n14573), .CK(clk), .Q(gray_img[1282]) );
  QDFFS gray_img_reg_10__1__2_ ( .D(n14572), .CK(clk), .Q(gray_img[1290]) );
  QDFFS gray_img_reg_10__2__2_ ( .D(n14571), .CK(clk), .Q(gray_img[1298]) );
  QDFFS gray_img_reg_10__3__2_ ( .D(n14570), .CK(clk), .Q(gray_img[1306]) );
  QDFFS gray_img_reg_10__4__2_ ( .D(n14569), .CK(clk), .Q(gray_img[1314]) );
  QDFFS gray_img_reg_10__5__2_ ( .D(n14568), .CK(clk), .Q(gray_img[1322]) );
  QDFFS gray_img_reg_10__6__2_ ( .D(n14567), .CK(clk), .Q(gray_img[1330]) );
  QDFFS gray_img_reg_10__7__2_ ( .D(n14566), .CK(clk), .Q(gray_img[1338]) );
  QDFFS gray_img_reg_10__8__2_ ( .D(n14565), .CK(clk), .Q(gray_img[1346]) );
  QDFFS gray_img_reg_10__9__2_ ( .D(n14564), .CK(clk), .Q(gray_img[1354]) );
  QDFFS gray_img_reg_10__10__2_ ( .D(n14563), .CK(clk), .Q(gray_img[1362]) );
  QDFFS gray_img_reg_10__11__2_ ( .D(n14562), .CK(clk), .Q(gray_img[1370]) );
  QDFFS gray_img_reg_10__12__2_ ( .D(n14561), .CK(clk), .Q(gray_img[1378]) );
  QDFFS gray_img_reg_10__13__2_ ( .D(n14560), .CK(clk), .Q(gray_img[1386]) );
  QDFFS gray_img_reg_10__14__2_ ( .D(n14559), .CK(clk), .Q(gray_img[1394]) );
  QDFFS gray_img_reg_10__15__2_ ( .D(n14558), .CK(clk), .Q(gray_img[1402]) );
  QDFFS gray_img_reg_11__0__2_ ( .D(n14557), .CK(clk), .Q(gray_img[1410]) );
  QDFFS gray_img_reg_11__1__2_ ( .D(n14556), .CK(clk), .Q(gray_img[1418]) );
  QDFFS gray_img_reg_11__2__2_ ( .D(n14555), .CK(clk), .Q(gray_img[1426]) );
  QDFFS gray_img_reg_11__3__2_ ( .D(n14554), .CK(clk), .Q(gray_img[1434]) );
  QDFFS gray_img_reg_11__4__2_ ( .D(n14553), .CK(clk), .Q(gray_img[1442]) );
  QDFFS gray_img_reg_11__5__2_ ( .D(n14552), .CK(clk), .Q(gray_img[1450]) );
  QDFFS gray_img_reg_11__6__2_ ( .D(n14551), .CK(clk), .Q(gray_img[1458]) );
  QDFFS gray_img_reg_11__7__2_ ( .D(n14550), .CK(clk), .Q(gray_img[1466]) );
  QDFFS gray_img_reg_11__8__2_ ( .D(n14549), .CK(clk), .Q(gray_img[1474]) );
  QDFFS gray_img_reg_11__9__2_ ( .D(n14548), .CK(clk), .Q(gray_img[1482]) );
  QDFFS gray_img_reg_11__10__2_ ( .D(n14547), .CK(clk), .Q(gray_img[1490]) );
  QDFFS gray_img_reg_11__11__2_ ( .D(n14546), .CK(clk), .Q(gray_img[1498]) );
  QDFFS gray_img_reg_11__12__2_ ( .D(n14545), .CK(clk), .Q(gray_img[1506]) );
  QDFFS gray_img_reg_11__13__2_ ( .D(n14544), .CK(clk), .Q(gray_img[1514]) );
  QDFFS gray_img_reg_11__14__2_ ( .D(n14543), .CK(clk), .Q(gray_img[1522]) );
  QDFFS gray_img_reg_11__15__2_ ( .D(n14542), .CK(clk), .Q(gray_img[1530]) );
  QDFFS gray_img_reg_12__0__2_ ( .D(n14541), .CK(clk), .Q(gray_img[1538]) );
  QDFFS gray_img_reg_12__1__2_ ( .D(n14540), .CK(clk), .Q(gray_img[1546]) );
  QDFFS gray_img_reg_12__2__2_ ( .D(n14539), .CK(clk), .Q(gray_img[1554]) );
  QDFFS gray_img_reg_12__3__2_ ( .D(n14538), .CK(clk), .Q(gray_img[1562]) );
  QDFFS gray_img_reg_12__4__2_ ( .D(n14537), .CK(clk), .Q(gray_img[1570]) );
  QDFFS gray_img_reg_12__5__2_ ( .D(n14536), .CK(clk), .Q(gray_img[1578]) );
  QDFFS gray_img_reg_12__6__2_ ( .D(n14535), .CK(clk), .Q(gray_img[1586]) );
  QDFFS gray_img_reg_12__7__2_ ( .D(n14534), .CK(clk), .Q(gray_img[1594]) );
  QDFFS gray_img_reg_12__8__2_ ( .D(n14533), .CK(clk), .Q(gray_img[1602]) );
  QDFFS gray_img_reg_12__9__2_ ( .D(n14532), .CK(clk), .Q(gray_img[1610]) );
  QDFFS gray_img_reg_12__10__2_ ( .D(n14531), .CK(clk), .Q(gray_img[1618]) );
  QDFFS gray_img_reg_12__11__2_ ( .D(n14530), .CK(clk), .Q(gray_img[1626]) );
  QDFFS gray_img_reg_12__12__2_ ( .D(n14529), .CK(clk), .Q(gray_img[1634]) );
  QDFFS gray_img_reg_12__13__2_ ( .D(n14528), .CK(clk), .Q(gray_img[1642]) );
  QDFFS gray_img_reg_12__14__2_ ( .D(n14527), .CK(clk), .Q(gray_img[1650]) );
  QDFFS gray_img_reg_12__15__2_ ( .D(n14526), .CK(clk), .Q(gray_img[1658]) );
  QDFFS gray_img_reg_13__0__2_ ( .D(n14525), .CK(clk), .Q(gray_img[1666]) );
  QDFFS gray_img_reg_13__1__2_ ( .D(n14524), .CK(clk), .Q(gray_img[1674]) );
  QDFFS gray_img_reg_13__2__2_ ( .D(n14523), .CK(clk), .Q(gray_img[1682]) );
  QDFFS gray_img_reg_13__3__2_ ( .D(n14522), .CK(clk), .Q(gray_img[1690]) );
  QDFFS gray_img_reg_13__4__2_ ( .D(n14521), .CK(clk), .Q(gray_img[1698]) );
  QDFFS gray_img_reg_13__5__2_ ( .D(n14520), .CK(clk), .Q(gray_img[1706]) );
  QDFFS gray_img_reg_13__6__2_ ( .D(n14519), .CK(clk), .Q(gray_img[1714]) );
  QDFFS gray_img_reg_13__7__2_ ( .D(n14518), .CK(clk), .Q(gray_img[1722]) );
  QDFFS gray_img_reg_13__8__2_ ( .D(n14517), .CK(clk), .Q(gray_img[1730]) );
  QDFFS gray_img_reg_13__9__2_ ( .D(n14516), .CK(clk), .Q(gray_img[1738]) );
  QDFFS gray_img_reg_13__10__2_ ( .D(n14515), .CK(clk), .Q(gray_img[1746]) );
  QDFFS gray_img_reg_13__11__2_ ( .D(n14514), .CK(clk), .Q(gray_img[1754]) );
  QDFFS gray_img_reg_13__12__2_ ( .D(n14513), .CK(clk), .Q(gray_img[1762]) );
  QDFFS gray_img_reg_13__13__2_ ( .D(n14512), .CK(clk), .Q(gray_img[1770]) );
  QDFFS gray_img_reg_13__14__2_ ( .D(n14511), .CK(clk), .Q(gray_img[1778]) );
  QDFFS gray_img_reg_13__15__2_ ( .D(n14510), .CK(clk), .Q(gray_img[1786]) );
  QDFFS gray_img_reg_14__0__2_ ( .D(n14509), .CK(clk), .Q(gray_img[1794]) );
  QDFFS gray_img_reg_14__1__2_ ( .D(n14508), .CK(clk), .Q(gray_img[1802]) );
  QDFFS gray_img_reg_14__2__2_ ( .D(n14507), .CK(clk), .Q(gray_img[1810]) );
  QDFFS gray_img_reg_14__3__2_ ( .D(n14506), .CK(clk), .Q(gray_img[1818]) );
  QDFFS gray_img_reg_14__4__2_ ( .D(n14505), .CK(clk), .Q(gray_img[1826]) );
  QDFFS gray_img_reg_14__5__2_ ( .D(n14504), .CK(clk), .Q(gray_img[1834]) );
  QDFFS gray_img_reg_14__6__2_ ( .D(n14503), .CK(clk), .Q(gray_img[1842]) );
  QDFFS gray_img_reg_14__7__2_ ( .D(n14502), .CK(clk), .Q(gray_img[1850]) );
  QDFFS gray_img_reg_14__8__2_ ( .D(n14501), .CK(clk), .Q(gray_img[1858]) );
  QDFFS gray_img_reg_14__9__2_ ( .D(n14500), .CK(clk), .Q(gray_img[1866]) );
  QDFFS gray_img_reg_14__10__2_ ( .D(n14499), .CK(clk), .Q(gray_img[1874]) );
  QDFFS gray_img_reg_14__11__2_ ( .D(n14498), .CK(clk), .Q(gray_img[1882]) );
  QDFFS gray_img_reg_14__12__2_ ( .D(n14497), .CK(clk), .Q(gray_img[1890]) );
  QDFFS gray_img_reg_14__13__2_ ( .D(n14496), .CK(clk), .Q(gray_img[1898]) );
  QDFFS gray_img_reg_14__14__2_ ( .D(n14495), .CK(clk), .Q(gray_img[1906]) );
  QDFFS gray_img_reg_14__15__2_ ( .D(n14494), .CK(clk), .Q(gray_img[1914]) );
  QDFFS gray_img_reg_15__0__2_ ( .D(n14493), .CK(clk), .Q(gray_img[1922]) );
  QDFFS gray_img_reg_15__1__2_ ( .D(n14492), .CK(clk), .Q(gray_img[1930]) );
  QDFFS gray_img_reg_15__2__2_ ( .D(n14491), .CK(clk), .Q(gray_img[1938]) );
  QDFFS gray_img_reg_15__3__2_ ( .D(n14490), .CK(clk), .Q(gray_img[1946]) );
  QDFFS gray_img_reg_15__4__2_ ( .D(n14489), .CK(clk), .Q(gray_img[1954]) );
  QDFFS gray_img_reg_15__5__2_ ( .D(n14488), .CK(clk), .Q(gray_img[1962]) );
  QDFFS gray_img_reg_15__6__2_ ( .D(n14487), .CK(clk), .Q(gray_img[1970]) );
  QDFFS gray_img_reg_15__8__2_ ( .D(n14485), .CK(clk), .Q(gray_img[1986]) );
  QDFFS gray_img_reg_15__9__2_ ( .D(n14484), .CK(clk), .Q(gray_img[1994]) );
  QDFFS gray_img_reg_15__10__2_ ( .D(n14483), .CK(clk), .Q(gray_img[2002]) );
  QDFFS gray_img_reg_15__11__2_ ( .D(n14482), .CK(clk), .Q(gray_img[2010]) );
  QDFFS gray_img_reg_15__12__2_ ( .D(n14481), .CK(clk), .Q(gray_img[2018]) );
  QDFFS gray_img_reg_15__13__2_ ( .D(n14480), .CK(clk), .Q(gray_img[2026]) );
  QDFFS gray_img_reg_15__14__2_ ( .D(n14479), .CK(clk), .Q(gray_img[2034]) );
  QDFFS gray_img_reg_15__15__2_ ( .D(n14478), .CK(clk), .Q(gray_img[2042]) );
  QDFFS gray_img_reg_5__5__2_ ( .D(n14470), .CK(clk), .Q(gray_img[682]) );
  QDFFS gray_img_reg_0__4__2_ ( .D(n14255), .CK(clk), .Q(gray_img[34]) );
  QDFFS gray_img_reg_0__5__2_ ( .D(n14246), .CK(clk), .Q(gray_img[42]) );
  QDFFS gray_img_reg_0__6__2_ ( .D(n14237), .CK(clk), .Q(gray_img[50]) );
  QDFFS gray_img_reg_0__7__2_ ( .D(n14228), .CK(clk), .Q(gray_img[58]) );
  QDFFS gray_img_reg_1__4__2_ ( .D(n14211), .CK(clk), .Q(gray_img[162]) );
  QDFFS gray_img_reg_1__5__2_ ( .D(n14202), .CK(clk), .Q(gray_img[170]) );
  QDFFS gray_img_reg_1__6__2_ ( .D(n14193), .CK(clk), .Q(gray_img[178]) );
  QDFFS gray_img_reg_1__7__2_ ( .D(n14184), .CK(clk), .Q(gray_img[186]) );
  QDFFS gray_img_reg_2__4__2_ ( .D(n14167), .CK(clk), .Q(gray_img[290]) );
  QDFFS gray_img_reg_2__5__2_ ( .D(n14158), .CK(clk), .Q(gray_img[298]) );
  QDFFS gray_img_reg_2__6__2_ ( .D(n14149), .CK(clk), .Q(gray_img[306]) );
  QDFFS gray_img_reg_2__7__2_ ( .D(n14140), .CK(clk), .Q(gray_img[314]) );
  QDFFS gray_img_reg_3__4__2_ ( .D(n14123), .CK(clk), .Q(gray_img[418]) );
  QDFFS gray_img_reg_3__5__2_ ( .D(n14114), .CK(clk), .Q(gray_img[426]) );
  QDFFS gray_img_reg_3__6__2_ ( .D(n14105), .CK(clk), .Q(gray_img[434]) );
  QDFFS gray_img_reg_3__7__2_ ( .D(n14096), .CK(clk), .Q(gray_img[442]) );
  QDFFS gray_img_reg_4__0__2_ ( .D(n14071), .CK(clk), .Q(gray_img[514]) );
  QDFFS gray_img_reg_4__1__2_ ( .D(n14062), .CK(clk), .Q(gray_img[522]) );
  QDFFS gray_img_reg_4__3__2_ ( .D(n14044), .CK(clk), .Q(gray_img[538]) );
  QDFFS gray_img_reg_4__4__2_ ( .D(n14035), .CK(clk), .Q(gray_img[546]) );
  QDFFS gray_img_reg_4__5__2_ ( .D(n14026), .CK(clk), .Q(gray_img[554]) );
  QDFFS gray_img_reg_4__6__2_ ( .D(n14017), .CK(clk), .Q(gray_img[562]) );
  QDFFS gray_img_reg_4__7__2_ ( .D(n14008), .CK(clk), .Q(gray_img[570]) );
  QDFFS gray_img_reg_5__0__2_ ( .D(n13983), .CK(clk), .Q(gray_img[642]) );
  QDFFS gray_img_reg_5__1__2_ ( .D(n13974), .CK(clk), .Q(gray_img[650]) );
  QDFFS gray_img_reg_5__2__2_ ( .D(n13965), .CK(clk), .Q(gray_img[658]) );
  QDFFS gray_img_reg_5__3__2_ ( .D(n13957), .CK(clk), .Q(gray_img[666]) );
  QDFFS gray_img_reg_5__4__2_ ( .D(n13949), .CK(clk), .Q(gray_img[674]) );
  QDFFS gray_img_reg_0__2__2_ ( .D(n13800), .CK(clk), .Q(gray_img[18]) );
  QDFFS gray_img_reg_0__3__2_ ( .D(n13790), .CK(clk), .Q(gray_img[26]) );
  QDFFS gray_img_reg_1__2__2_ ( .D(n13770), .CK(clk), .Q(gray_img[146]) );
  QDFFS gray_img_reg_1__3__2_ ( .D(n13760), .CK(clk), .Q(gray_img[154]) );
  QDFFS gray_img_reg_0__1__2_ ( .D(n13752), .CK(clk), .Q(gray_img[10]) );
  QDFFS gray_img_reg_2__0__2_ ( .D(n13734), .CK(clk), .Q(gray_img[258]) );
  QDFFS gray_img_reg_2__1__2_ ( .D(n13705), .CK(clk), .Q(gray_img[266]) );
  QDFFS gray_img_reg_2__2__2_ ( .D(n13679), .CK(clk), .Q(gray_img[274]) );
  QDFFS gray_img_reg_5__6__2_ ( .D(n13673), .CK(clk), .Q(gray_img[690]) );
  QDFFS gray_img_reg_5__7__2_ ( .D(n13672), .CK(clk), .Q(gray_img[698]) );
  QDFFS gray_img_reg_2__3__2_ ( .D(n14670), .CK(clk), .Q(gray_img[282]) );
  QDFFS gray_img_reg_6__0__2_ ( .D(n13671), .CK(clk), .Q(gray_img[770]) );
  QDFFS gray_img_reg_6__1__2_ ( .D(n13670), .CK(clk), .Q(gray_img[778]) );
  QDFFS gray_img_reg_6__2__2_ ( .D(n13669), .CK(clk), .Q(gray_img[786]) );
  QDFFS gray_img_reg_6__3__2_ ( .D(n13668), .CK(clk), .Q(gray_img[794]) );
  QDFFS gray_img_reg_6__4__2_ ( .D(n13667), .CK(clk), .Q(gray_img[802]) );
  QDFFS gray_img_reg_6__5__2_ ( .D(n13666), .CK(clk), .Q(gray_img[810]) );
  QDFFS gray_img_reg_6__6__2_ ( .D(n13665), .CK(clk), .Q(gray_img[818]) );
  QDFFS gray_img_reg_6__7__2_ ( .D(n13664), .CK(clk), .Q(gray_img[826]) );
  QDFFS gray_img_reg_7__0__2_ ( .D(n13663), .CK(clk), .Q(gray_img[898]) );
  QDFFS gray_img_reg_7__1__2_ ( .D(n13662), .CK(clk), .Q(gray_img[906]) );
  QDFFS gray_img_reg_3__0__2_ ( .D(n14474), .CK(clk), .Q(gray_img[386]) );
  QDFFS gray_img_reg_7__2__2_ ( .D(n13661), .CK(clk), .Q(gray_img[914]) );
  QDFFS gray_img_reg_7__3__2_ ( .D(n13660), .CK(clk), .Q(gray_img[922]) );
  QDFFS gray_img_reg_3__1__2_ ( .D(n14473), .CK(clk), .Q(gray_img[394]) );
  QDFFS gray_img_reg_1__0__2_ ( .D(n14476), .CK(clk), .Q(gray_img[130]) );
  QDFFS gray_img_reg_7__4__2_ ( .D(n13659), .CK(clk), .Q(gray_img[930]) );
  QDFFS gray_img_reg_7__5__2_ ( .D(n13658), .CK(clk), .Q(gray_img[938]) );
  QDFFS gray_img_reg_3__2__2_ ( .D(n14472), .CK(clk), .Q(gray_img[402]) );
  QDFFS gray_img_reg_7__6__2_ ( .D(n13657), .CK(clk), .Q(gray_img[946]) );
  QDFFS gray_img_reg_7__7__2_ ( .D(n13656), .CK(clk), .Q(gray_img[954]) );
  QDFFS gray_img_reg_3__3__2_ ( .D(n14471), .CK(clk), .Q(gray_img[410]) );
  QDFFS gray_img_reg_1__1__2_ ( .D(n14475), .CK(clk), .Q(gray_img[138]) );
  QDFFS mem_data_out_reg_shift_0_reg_0__1_ ( .D(n15814), .CK(clk), .Q(
        mem_data_out_reg_shift_0[1]) );
  QDFFS mem_data_out_reg_shift_0_reg_1__1_ ( .D(mem_data_out_reg_shift_0[1]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[9]) );
  QDFFS mem_data_out_reg_shift_0_reg_2__1_ ( .D(mem_data_out_reg_shift_0[9]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[17]) );
  QDFFS mem_data_out_reg_shift_0_reg_3__1_ ( .D(mem_data_out_reg_shift_0[17]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[25]) );
  QDFFS mem_data_out_reg_shift_0_reg_4__1_ ( .D(mem_data_out_reg_shift_0[25]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[33]) );
  QDFFS mem_data_out_reg_shift_0_reg_5__1_ ( .D(mem_data_out_reg_shift_0[33]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[41]) );
  QDFFS mem_data_out_reg_shift_0_reg_6__1_ ( .D(mem_data_out_reg_shift_0[41]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[49]) );
  QDFFS mem_data_out_reg_shift_0_reg_7__1_ ( .D(mem_data_out_reg_shift_0[49]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[57]) );
  QDFFS mem_data_out_reg_shift_0_reg_8__1_ ( .D(mem_data_out_reg_shift_0[57]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[65]) );
  QDFFS mem_data_out_reg_shift_0_reg_9__1_ ( .D(mem_data_out_reg_shift_0[65]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[73]) );
  QDFFS mem_data_out_reg_shift_0_reg_10__1_ ( .D(mem_data_out_reg_shift_0[73]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[81]) );
  QDFFS mem_data_out_reg_shift_0_reg_11__1_ ( .D(mem_data_out_reg_shift_0[81]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[89]) );
  QDFFS mem_data_out_reg_shift_0_reg_12__1_ ( .D(mem_data_out_reg_shift_0[89]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[97]) );
  QDFFS mem_data_out_reg_shift_0_reg_13__1_ ( .D(mem_data_out_reg_shift_0[97]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[105]) );
  QDFFS mem_data_out_reg_shift_0_reg_14__1_ ( .D(mem_data_out_reg_shift_0[105]), .CK(clk), .Q(mem_data_out_reg_shift_0[113]) );
  QDFFS mem_data_out_reg_shift_0_reg_15__1_ ( .D(mem_data_out_reg_shift_0[113]), .CK(clk), .Q(mem_data_out_reg_shift_0[121]) );
  QDFFS mem_data_out_reg_shift_1_reg_0__1_ ( .D(n15831), .CK(clk), .Q(
        mem_data_out_reg_shift_1[1]) );
  QDFFS mem_data_out_reg_shift_1_reg_1__1_ ( .D(mem_data_out_reg_shift_1[1]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[9]) );
  QDFFS mem_data_out_reg_shift_1_reg_3__1_ ( .D(mem_data_out_reg_shift_1[17]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[25]) );
  QDFFS mem_data_out_reg_shift_1_reg_4__1_ ( .D(mem_data_out_reg_shift_1[25]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[33]) );
  QDFFS mem_data_out_reg_shift_1_reg_5__1_ ( .D(mem_data_out_reg_shift_1[33]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[41]) );
  QDFFS mem_data_out_reg_shift_1_reg_6__1_ ( .D(mem_data_out_reg_shift_1[41]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[49]) );
  QDFFS mem_data_out_reg_shift_1_reg_7__1_ ( .D(mem_data_out_reg_shift_1[49]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[57]) );
  QDFFS mem_data_out_reg_shift_1_reg_8__1_ ( .D(mem_data_out_reg_shift_1[57]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[65]) );
  QDFFS mem_data_out_reg_shift_1_reg_9__1_ ( .D(mem_data_out_reg_shift_1[65]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[73]) );
  QDFFS mem_data_out_reg_shift_1_reg_10__1_ ( .D(mem_data_out_reg_shift_1[73]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[81]) );
  QDFFS mem_data_out_reg_shift_1_reg_11__1_ ( .D(mem_data_out_reg_shift_1[81]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[89]) );
  QDFFS mem_data_out_reg_shift_1_reg_12__1_ ( .D(mem_data_out_reg_shift_1[89]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[97]) );
  QDFFS mem_data_out_reg_shift_1_reg_13__1_ ( .D(mem_data_out_reg_shift_1[97]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[105]) );
  QDFFS mem_data_out_reg_shift_1_reg_14__1_ ( .D(mem_data_out_reg_shift_1[105]), .CK(clk), .Q(mem_data_out_reg_shift_1[113]) );
  QDFFS mem_data_out_reg_shift_1_reg_15__1_ ( .D(mem_data_out_reg_shift_1[113]), .CK(clk), .Q(mem_data_out_reg_shift_1[121]) );
  QDFFS mem_data_out_reg_shift_2_reg_0__1_ ( .D(n15839), .CK(clk), .Q(
        mem_data_out_reg_shift_2[1]) );
  QDFFS mem_data_out_reg_shift_2_reg_1__1_ ( .D(mem_data_out_reg_shift_2[1]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[9]) );
  QDFFS mem_data_out_reg_shift_2_reg_2__1_ ( .D(mem_data_out_reg_shift_2[9]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[17]) );
  QDFFS mem_data_out_reg_shift_2_reg_3__1_ ( .D(mem_data_out_reg_shift_2[17]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[25]) );
  QDFFS medfilt_out_reg_reg_1_ ( .D(n15858), .CK(clk), .Q(medfilt_out_reg[1])
         );
  QDFFS gray_img_reg_0__13__1_ ( .D(n14463), .CK(clk), .Q(gray_img[105]) );
  QDFFS gray_img_reg_1__9__1_ ( .D(n14459), .CK(clk), .Q(gray_img[201]) );
  QDFFS gray_img_reg_1__13__1_ ( .D(n14455), .CK(clk), .Q(gray_img[233]) );
  QDFFS gray_img_reg_2__8__1_ ( .D(n14452), .CK(clk), .Q(gray_img[321]) );
  QDFFS gray_img_reg_2__9__1_ ( .D(n14451), .CK(clk), .Q(gray_img[329]) );
  QDFFS gray_img_reg_2__15__1_ ( .D(n14445), .CK(clk), .Q(gray_img[377]) );
  QDFFS gray_img_reg_3__13__1_ ( .D(n14439), .CK(clk), .Q(gray_img[489]) );
  QDFFS gray_img_reg_4__9__1_ ( .D(n14435), .CK(clk), .Q(gray_img[585]) );
  QDFFS gray_img_reg_4__12__1_ ( .D(n14432), .CK(clk), .Q(gray_img[609]) );
  QDFFS gray_img_reg_5__12__1_ ( .D(n14424), .CK(clk), .Q(gray_img[737]) );
  QDFFS gray_img_reg_5__13__1_ ( .D(n14423), .CK(clk), .Q(gray_img[745]) );
  QDFFS gray_img_reg_6__9__1_ ( .D(n14419), .CK(clk), .Q(gray_img[841]) );
  QDFFS gray_img_reg_6__13__1_ ( .D(n14415), .CK(clk), .Q(gray_img[873]) );
  QDFFS gray_img_reg_6__14__1_ ( .D(n14414), .CK(clk), .Q(gray_img[881]) );
  QDFFS gray_img_reg_7__8__1_ ( .D(n14412), .CK(clk), .Q(gray_img[961]) );
  QDFFS gray_img_reg_7__13__1_ ( .D(n14407), .CK(clk), .Q(gray_img[1001]) );
  QDFFS gray_img_reg_7__14__1_ ( .D(n14406), .CK(clk), .Q(gray_img[1009]) );
  QDFFS gray_img_reg_8__0__1_ ( .D(n14404), .CK(clk), .Q(gray_img[1025]) );
  QDFFS gray_img_reg_8__4__1_ ( .D(n14400), .CK(clk), .Q(gray_img[1057]) );
  QDFFS gray_img_reg_8__6__1_ ( .D(n14398), .CK(clk), .Q(gray_img[1073]) );
  QDFFS gray_img_reg_8__7__1_ ( .D(n14397), .CK(clk), .Q(gray_img[1081]) );
  QDFFS gray_img_reg_8__9__1_ ( .D(n14395), .CK(clk), .Q(gray_img[1097]) );
  QDFFS gray_img_reg_8__11__1_ ( .D(n14393), .CK(clk), .Q(gray_img[1113]) );
  QDFFS gray_img_reg_8__12__1_ ( .D(n14392), .CK(clk), .Q(gray_img[1121]) );
  QDFFS gray_img_reg_9__9__1_ ( .D(n14379), .CK(clk), .Q(gray_img[1225]) );
  QDFFS gray_img_reg_9__10__1_ ( .D(n14378), .CK(clk), .Q(gray_img[1233]) );
  QDFFS gray_img_reg_9__11__1_ ( .D(n14377), .CK(clk), .Q(gray_img[1241]) );
  QDFFS gray_img_reg_9__14__1_ ( .D(n14374), .CK(clk), .Q(gray_img[1265]) );
  QDFFS gray_img_reg_10__2__1_ ( .D(n14370), .CK(clk), .Q(gray_img[1297]) );
  QDFFS gray_img_reg_10__6__1_ ( .D(n14366), .CK(clk), .Q(gray_img[1329]) );
  QDFFS gray_img_reg_10__8__1_ ( .D(n14364), .CK(clk), .Q(gray_img[1345]) );
  QDFFS gray_img_reg_10__9__1_ ( .D(n14363), .CK(clk), .Q(gray_img[1353]) );
  QDFFS gray_img_reg_10__12__1_ ( .D(n14360), .CK(clk), .Q(gray_img[1377]) );
  QDFFS gray_img_reg_10__13__1_ ( .D(n14359), .CK(clk), .Q(gray_img[1385]) );
  QDFFS gray_img_reg_10__14__1_ ( .D(n14358), .CK(clk), .Q(gray_img[1393]) );
  QDFFS gray_img_reg_10__15__1_ ( .D(n14357), .CK(clk), .Q(gray_img[1401]) );
  QDFFS gray_img_reg_11__1__1_ ( .D(n14355), .CK(clk), .Q(gray_img[1417]) );
  QDFFS gray_img_reg_11__2__1_ ( .D(n14354), .CK(clk), .Q(gray_img[1425]) );
  QDFFS gray_img_reg_11__3__1_ ( .D(n14353), .CK(clk), .Q(gray_img[1433]) );
  QDFFS gray_img_reg_11__6__1_ ( .D(n14350), .CK(clk), .Q(gray_img[1457]) );
  QDFFS gray_img_reg_11__11__1_ ( .D(n14345), .CK(clk), .Q(gray_img[1497]) );
  QDFFS gray_img_reg_11__12__1_ ( .D(n14344), .CK(clk), .Q(gray_img[1505]) );
  QDFFS gray_img_reg_11__14__1_ ( .D(n14342), .CK(clk), .Q(gray_img[1521]) );
  QDFFS gray_img_reg_12__1__1_ ( .D(n14339), .CK(clk), .Q(gray_img[1545]) );
  QDFFS gray_img_reg_12__2__1_ ( .D(n14338), .CK(clk), .Q(gray_img[1553]) );
  QDFFS gray_img_reg_12__3__1_ ( .D(n14337), .CK(clk), .Q(gray_img[1561]) );
  QDFFS gray_img_reg_12__4__1_ ( .D(n14336), .CK(clk), .Q(gray_img[1569]) );
  QDFFS gray_img_reg_12__5__1_ ( .D(n14335), .CK(clk), .Q(gray_img[1577]) );
  QDFFS gray_img_reg_12__6__1_ ( .D(n14334), .CK(clk), .Q(gray_img[1585]) );
  QDFFS gray_img_reg_12__7__1_ ( .D(n14333), .CK(clk), .Q(gray_img[1593]) );
  QDFFS gray_img_reg_12__10__1_ ( .D(n14330), .CK(clk), .Q(gray_img[1617]) );
  QDFFS gray_img_reg_12__11__1_ ( .D(n14329), .CK(clk), .Q(gray_img[1625]) );
  QDFFS gray_img_reg_12__14__1_ ( .D(n14326), .CK(clk), .Q(gray_img[1649]) );
  QDFFS gray_img_reg_12__15__1_ ( .D(n14325), .CK(clk), .Q(gray_img[1657]) );
  QDFFS gray_img_reg_13__3__1_ ( .D(n14321), .CK(clk), .Q(gray_img[1689]) );
  QDFFS gray_img_reg_13__8__1_ ( .D(n14316), .CK(clk), .Q(gray_img[1729]) );
  QDFFS gray_img_reg_13__9__1_ ( .D(n14315), .CK(clk), .Q(gray_img[1737]) );
  QDFFS gray_img_reg_13__10__1_ ( .D(n14314), .CK(clk), .Q(gray_img[1745]) );
  QDFFS gray_img_reg_13__11__1_ ( .D(n14313), .CK(clk), .Q(gray_img[1753]) );
  QDFFS gray_img_reg_13__13__1_ ( .D(n14311), .CK(clk), .Q(gray_img[1769]) );
  QDFFS gray_img_reg_14__1__1_ ( .D(n14307), .CK(clk), .Q(gray_img[1801]) );
  QDFFS gray_img_reg_14__4__1_ ( .D(n14304), .CK(clk), .Q(gray_img[1825]) );
  QDFFS gray_img_reg_14__5__1_ ( .D(n14303), .CK(clk), .Q(gray_img[1833]) );
  QDFFS gray_img_reg_14__9__1_ ( .D(n14299), .CK(clk), .Q(gray_img[1865]) );
  QDFFS gray_img_reg_14__10__1_ ( .D(n14298), .CK(clk), .Q(gray_img[1873]) );
  QDFFS gray_img_reg_14__11__1_ ( .D(n14297), .CK(clk), .Q(gray_img[1881]) );
  QDFFS gray_img_reg_14__12__1_ ( .D(n14296), .CK(clk), .Q(gray_img[1889]) );
  QDFFS gray_img_reg_14__13__1_ ( .D(n14295), .CK(clk), .Q(gray_img[1897]) );
  QDFFS gray_img_reg_14__14__1_ ( .D(n14294), .CK(clk), .Q(gray_img[1905]) );
  QDFFS gray_img_reg_15__1__1_ ( .D(n14291), .CK(clk), .Q(gray_img[1929]) );
  QDFFS gray_img_reg_15__4__1_ ( .D(n14288), .CK(clk), .Q(gray_img[1953]) );
  QDFFS gray_img_reg_15__5__1_ ( .D(n14287), .CK(clk), .Q(gray_img[1961]) );
  QDFFS gray_img_reg_15__9__1_ ( .D(n14283), .CK(clk), .Q(gray_img[1993]) );
  QDFFS gray_img_reg_15__10__1_ ( .D(n14282), .CK(clk), .Q(gray_img[2001]) );
  QDFFS gray_img_reg_15__11__1_ ( .D(n14281), .CK(clk), .Q(gray_img[2009]) );
  QDFFS gray_img_reg_5__3__1_ ( .D(n14268), .CK(clk), .Q(gray_img[665]) );
  QDFFS gray_img_reg_0__4__1_ ( .D(n14256), .CK(clk), .Q(gray_img[33]) );
  QDFFS gray_img_reg_0__7__1_ ( .D(n14229), .CK(clk), .Q(gray_img[57]) );
  QDFFS gray_img_reg_1__5__1_ ( .D(n14203), .CK(clk), .Q(gray_img[169]) );
  QDFFS gray_img_reg_1__6__1_ ( .D(n14194), .CK(clk), .Q(gray_img[177]) );
  QDFFS gray_img_reg_2__4__1_ ( .D(n14168), .CK(clk), .Q(gray_img[289]) );
  QDFFS gray_img_reg_3__4__1_ ( .D(n14124), .CK(clk), .Q(gray_img[417]) );
  QDFFS gray_img_reg_3__6__1_ ( .D(n14106), .CK(clk), .Q(gray_img[433]) );
  QDFFS gray_img_reg_4__1__1_ ( .D(n14063), .CK(clk), .Q(gray_img[521]) );
  QDFFS gray_img_reg_4__3__1_ ( .D(n14045), .CK(clk), .Q(gray_img[537]) );
  QDFFS gray_img_reg_5__1__1_ ( .D(n13975), .CK(clk), .Q(gray_img[649]) );
  QDFFS gray_img_reg_0__3__1_ ( .D(n13791), .CK(clk), .Q(gray_img[25]) );
  QDFFS gray_img_reg_1__2__1_ ( .D(n13771), .CK(clk), .Q(gray_img[145]) );
  QDFFS gray_img_reg_1__3__1_ ( .D(n13761), .CK(clk), .Q(gray_img[153]) );
  QDFFS gray_img_reg_0__1__1_ ( .D(n13753), .CK(clk), .Q(gray_img[9]) );
  QDFFS gray_img_reg_2__1__1_ ( .D(n13706), .CK(clk), .Q(gray_img[265]) );
  QDFFS gray_img_reg_5__5__1_ ( .D(n13698), .CK(clk), .Q(gray_img[681]) );
  QDFFS gray_img_reg_5__7__1_ ( .D(n13696), .CK(clk), .Q(gray_img[697]) );
  QDFFS gray_img_reg_2__3__1_ ( .D(n14273), .CK(clk), .Q(gray_img[281]) );
  QDFFS gray_img_reg_6__0__1_ ( .D(n13695), .CK(clk), .Q(gray_img[769]) );
  QDFFS gray_img_reg_6__1__1_ ( .D(n13694), .CK(clk), .Q(gray_img[777]) );
  QDFFS gray_img_reg_6__2__1_ ( .D(n13693), .CK(clk), .Q(gray_img[785]) );
  QDFFS gray_img_reg_6__3__1_ ( .D(n13692), .CK(clk), .Q(gray_img[793]) );
  QDFFS gray_img_reg_6__4__1_ ( .D(n13691), .CK(clk), .Q(gray_img[801]) );
  QDFFS gray_img_reg_6__5__1_ ( .D(n13690), .CK(clk), .Q(gray_img[809]) );
  QDFFS gray_img_reg_6__6__1_ ( .D(n13689), .CK(clk), .Q(gray_img[817]) );
  QDFFS gray_img_reg_6__7__1_ ( .D(n13688), .CK(clk), .Q(gray_img[825]) );
  QDFFS gray_img_reg_1__0__1_ ( .D(n14275), .CK(clk), .Q(gray_img[129]) );
  QDFFS gray_img_reg_7__4__1_ ( .D(n13683), .CK(clk), .Q(gray_img[929]) );
  QDFFS gray_img_reg_7__6__1_ ( .D(n13681), .CK(clk), .Q(gray_img[945]) );
  QDFFS gray_img_reg_7__7__1_ ( .D(n13680), .CK(clk), .Q(gray_img[953]) );
  QDFFS gray_img_reg_1__1__1_ ( .D(n14274), .CK(clk), .Q(gray_img[137]) );
  QDFFS gray_img_reg_0__0__0_ ( .D(n13811), .CK(clk), .Q(gray_img[0]) );
  QDFFS mem_data_out_reg_shift_0_reg_0__0_ ( .D(n15815), .CK(clk), .Q(
        mem_data_out_reg_shift_0[0]) );
  QDFFS mem_data_out_reg_shift_0_reg_1__0_ ( .D(mem_data_out_reg_shift_0[0]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[8]) );
  QDFFS mem_data_out_reg_shift_0_reg_2__0_ ( .D(mem_data_out_reg_shift_0[8]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[16]) );
  QDFFS mem_data_out_reg_shift_0_reg_3__0_ ( .D(mem_data_out_reg_shift_0[16]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[24]) );
  QDFFS mem_data_out_reg_shift_0_reg_4__0_ ( .D(mem_data_out_reg_shift_0[24]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[32]) );
  QDFFS mem_data_out_reg_shift_0_reg_5__0_ ( .D(mem_data_out_reg_shift_0[32]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[40]) );
  QDFFS mem_data_out_reg_shift_0_reg_6__0_ ( .D(mem_data_out_reg_shift_0[40]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[48]) );
  QDFFS mem_data_out_reg_shift_0_reg_7__0_ ( .D(mem_data_out_reg_shift_0[48]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[56]) );
  QDFFS mem_data_out_reg_shift_0_reg_8__0_ ( .D(mem_data_out_reg_shift_0[56]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[64]) );
  QDFFS mem_data_out_reg_shift_0_reg_9__0_ ( .D(mem_data_out_reg_shift_0[64]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[72]) );
  QDFFS mem_data_out_reg_shift_0_reg_10__0_ ( .D(mem_data_out_reg_shift_0[72]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[80]) );
  QDFFS mem_data_out_reg_shift_0_reg_11__0_ ( .D(mem_data_out_reg_shift_0[80]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[88]) );
  QDFFS mem_data_out_reg_shift_0_reg_12__0_ ( .D(mem_data_out_reg_shift_0[88]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[96]) );
  QDFFS mem_data_out_reg_shift_0_reg_13__0_ ( .D(mem_data_out_reg_shift_0[96]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[104]) );
  QDFFS mem_data_out_reg_shift_0_reg_14__0_ ( .D(mem_data_out_reg_shift_0[104]), .CK(clk), .Q(mem_data_out_reg_shift_0[112]) );
  QDFFS mem_data_out_reg_shift_0_reg_15__0_ ( .D(mem_data_out_reg_shift_0[112]), .CK(clk), .Q(mem_data_out_reg_shift_0[120]) );
  QDFFS mem_data_out_reg_shift_1_reg_0__0_ ( .D(n15832), .CK(clk), .Q(
        mem_data_out_reg_shift_1[0]) );
  QDFFS mem_data_out_reg_shift_1_reg_1__0_ ( .D(mem_data_out_reg_shift_1[0]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[8]) );
  QDFFS mem_data_out_reg_shift_1_reg_3__0_ ( .D(mem_data_out_reg_shift_1[16]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[24]) );
  QDFFS mem_data_out_reg_shift_1_reg_4__0_ ( .D(mem_data_out_reg_shift_1[24]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[32]) );
  QDFFS mem_data_out_reg_shift_1_reg_5__0_ ( .D(mem_data_out_reg_shift_1[32]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[40]) );
  QDFFS mem_data_out_reg_shift_1_reg_6__0_ ( .D(mem_data_out_reg_shift_1[40]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[48]) );
  QDFFS mem_data_out_reg_shift_1_reg_7__0_ ( .D(mem_data_out_reg_shift_1[48]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[56]) );
  QDFFS mem_data_out_reg_shift_1_reg_8__0_ ( .D(mem_data_out_reg_shift_1[56]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[64]) );
  QDFFS mem_data_out_reg_shift_1_reg_9__0_ ( .D(mem_data_out_reg_shift_1[64]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[72]) );
  QDFFS mem_data_out_reg_shift_1_reg_10__0_ ( .D(mem_data_out_reg_shift_1[72]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[80]) );
  QDFFS mem_data_out_reg_shift_1_reg_11__0_ ( .D(mem_data_out_reg_shift_1[80]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[88]) );
  QDFFS mem_data_out_reg_shift_1_reg_12__0_ ( .D(mem_data_out_reg_shift_1[88]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[96]) );
  QDFFS mem_data_out_reg_shift_1_reg_13__0_ ( .D(mem_data_out_reg_shift_1[96]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[104]) );
  QDFFS mem_data_out_reg_shift_1_reg_14__0_ ( .D(mem_data_out_reg_shift_1[104]), .CK(clk), .Q(mem_data_out_reg_shift_1[112]) );
  QDFFS mem_data_out_reg_shift_1_reg_15__0_ ( .D(mem_data_out_reg_shift_1[112]), .CK(clk), .Q(mem_data_out_reg_shift_1[120]) );
  QDFFS mem_data_out_reg_shift_2_reg_0__0_ ( .D(n15840), .CK(clk), .Q(
        mem_data_out_reg_shift_2[0]) );
  QDFFS mem_data_out_reg_shift_2_reg_1__0_ ( .D(mem_data_out_reg_shift_2[0]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[8]) );
  QDFFS mem_data_out_reg_shift_2_reg_2__0_ ( .D(mem_data_out_reg_shift_2[8]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[16]) );
  QDFFS mem_data_out_reg_shift_2_reg_3__0_ ( .D(mem_data_out_reg_shift_2[16]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[24]) );
  QDFFS medfilt_out_reg_reg_0_ ( .D(n15857), .CK(clk), .Q(medfilt_out_reg[0])
         );
  QDFFS gray_img_reg_0__12__0_ ( .D(n14262), .CK(clk), .Q(gray_img[96]) );
  QDFFS gray_img_reg_0__13__0_ ( .D(n14261), .CK(clk), .Q(gray_img[104]) );
  QDFFS gray_img_reg_0__15__0_ ( .D(n14259), .CK(clk), .Q(gray_img[120]) );
  QDFFS gray_img_reg_1__8__0_ ( .D(n14258), .CK(clk), .Q(gray_img[192]) );
  QDFFS gray_img_reg_1__9__0_ ( .D(n14257), .CK(clk), .Q(gray_img[200]) );
  QDFFS gray_img_reg_1__10__0_ ( .D(n14249), .CK(clk), .Q(gray_img[208]) );
  QDFFS gray_img_reg_1__11__0_ ( .D(n14248), .CK(clk), .Q(gray_img[216]) );
  QDFFS gray_img_reg_1__12__0_ ( .D(n14240), .CK(clk), .Q(gray_img[224]) );
  QDFFS gray_img_reg_1__13__0_ ( .D(n14239), .CK(clk), .Q(gray_img[232]) );
  QDFFS gray_img_reg_1__14__0_ ( .D(n14231), .CK(clk), .Q(gray_img[240]) );
  QDFFS gray_img_reg_1__15__0_ ( .D(n14230), .CK(clk), .Q(gray_img[248]) );
  QDFFS gray_img_reg_2__8__0_ ( .D(n14222), .CK(clk), .Q(gray_img[320]) );
  QDFFS gray_img_reg_2__9__0_ ( .D(n14221), .CK(clk), .Q(gray_img[328]) );
  QDFFS gray_img_reg_2__12__0_ ( .D(n14218), .CK(clk), .Q(gray_img[352]) );
  QDFFS gray_img_reg_2__13__0_ ( .D(n14217), .CK(clk), .Q(gray_img[360]) );
  QDFFS gray_img_reg_2__14__0_ ( .D(n14216), .CK(clk), .Q(gray_img[368]) );
  QDFFS gray_img_reg_2__15__0_ ( .D(n14215), .CK(clk), .Q(gray_img[376]) );
  QDFFS gray_img_reg_3__8__0_ ( .D(n14214), .CK(clk), .Q(gray_img[448]) );
  QDFFS gray_img_reg_3__9__0_ ( .D(n14213), .CK(clk), .Q(gray_img[456]) );
  QDFFS gray_img_reg_3__10__0_ ( .D(n14205), .CK(clk), .Q(gray_img[464]) );
  QDFFS gray_img_reg_3__11__0_ ( .D(n14204), .CK(clk), .Q(gray_img[472]) );
  QDFFS gray_img_reg_3__12__0_ ( .D(n14196), .CK(clk), .Q(gray_img[480]) );
  QDFFS gray_img_reg_3__14__0_ ( .D(n14187), .CK(clk), .Q(gray_img[496]) );
  QDFFS gray_img_reg_3__15__0_ ( .D(n14186), .CK(clk), .Q(gray_img[504]) );
  QDFFS gray_img_reg_4__8__0_ ( .D(n14178), .CK(clk), .Q(gray_img[576]) );
  QDFFS gray_img_reg_4__9__0_ ( .D(n14177), .CK(clk), .Q(gray_img[584]) );
  QDFFS gray_img_reg_4__10__0_ ( .D(n14176), .CK(clk), .Q(gray_img[592]) );
  QDFFS gray_img_reg_4__11__0_ ( .D(n14175), .CK(clk), .Q(gray_img[600]) );
  QDFFS gray_img_reg_4__12__0_ ( .D(n14174), .CK(clk), .Q(gray_img[608]) );
  QDFFS gray_img_reg_4__13__0_ ( .D(n14173), .CK(clk), .Q(gray_img[616]) );
  QDFFS gray_img_reg_4__14__0_ ( .D(n14172), .CK(clk), .Q(gray_img[624]) );
  QDFFS gray_img_reg_4__15__0_ ( .D(n14171), .CK(clk), .Q(gray_img[632]) );
  QDFFS gray_img_reg_5__8__0_ ( .D(n14170), .CK(clk), .Q(gray_img[704]) );
  QDFFS gray_img_reg_5__9__0_ ( .D(n14169), .CK(clk), .Q(gray_img[712]) );
  QDFFS gray_img_reg_5__11__0_ ( .D(n14160), .CK(clk), .Q(gray_img[728]) );
  QDFFS gray_img_reg_5__12__0_ ( .D(n14152), .CK(clk), .Q(gray_img[736]) );
  QDFFS gray_img_reg_5__13__0_ ( .D(n14151), .CK(clk), .Q(gray_img[744]) );
  QDFFS gray_img_reg_5__14__0_ ( .D(n14143), .CK(clk), .Q(gray_img[752]) );
  QDFFS gray_img_reg_5__15__0_ ( .D(n14142), .CK(clk), .Q(gray_img[760]) );
  QDFFS gray_img_reg_6__8__0_ ( .D(n14134), .CK(clk), .Q(gray_img[832]) );
  QDFFS gray_img_reg_6__9__0_ ( .D(n14133), .CK(clk), .Q(gray_img[840]) );
  QDFFS gray_img_reg_6__10__0_ ( .D(n14132), .CK(clk), .Q(gray_img[848]) );
  QDFFS gray_img_reg_6__11__0_ ( .D(n14131), .CK(clk), .Q(gray_img[856]) );
  QDFFS gray_img_reg_6__12__0_ ( .D(n14130), .CK(clk), .Q(gray_img[864]) );
  QDFFS gray_img_reg_6__13__0_ ( .D(n14129), .CK(clk), .Q(gray_img[872]) );
  QDFFS gray_img_reg_6__14__0_ ( .D(n14128), .CK(clk), .Q(gray_img[880]) );
  QDFFS gray_img_reg_6__15__0_ ( .D(n14127), .CK(clk), .Q(gray_img[888]) );
  QDFFS gray_img_reg_7__9__0_ ( .D(n14125), .CK(clk), .Q(gray_img[968]) );
  QDFFS gray_img_reg_7__12__0_ ( .D(n14108), .CK(clk), .Q(gray_img[992]) );
  QDFFS gray_img_reg_7__13__0_ ( .D(n14107), .CK(clk), .Q(gray_img[1000]) );
  QDFFS gray_img_reg_7__14__0_ ( .D(n14099), .CK(clk), .Q(gray_img[1008]) );
  QDFFS gray_img_reg_7__15__0_ ( .D(n14098), .CK(clk), .Q(gray_img[1016]) );
  QDFFS gray_img_reg_8__0__0_ ( .D(n14090), .CK(clk), .Q(gray_img[1024]) );
  QDFFS gray_img_reg_8__1__0_ ( .D(n14089), .CK(clk), .Q(gray_img[1032]) );
  QDFFS gray_img_reg_8__4__0_ ( .D(n14086), .CK(clk), .Q(gray_img[1056]) );
  QDFFS gray_img_reg_8__6__0_ ( .D(n14084), .CK(clk), .Q(gray_img[1072]) );
  QDFFS gray_img_reg_8__9__0_ ( .D(n14081), .CK(clk), .Q(gray_img[1096]) );
  QDFFS gray_img_reg_8__10__0_ ( .D(n14080), .CK(clk), .Q(gray_img[1104]) );
  QDFFS gray_img_reg_8__11__0_ ( .D(n14079), .CK(clk), .Q(gray_img[1112]) );
  QDFFS gray_img_reg_8__12__0_ ( .D(n14078), .CK(clk), .Q(gray_img[1120]) );
  QDFFS gray_img_reg_8__13__0_ ( .D(n14077), .CK(clk), .Q(gray_img[1128]) );
  QDFFS gray_img_reg_8__14__0_ ( .D(n14076), .CK(clk), .Q(gray_img[1136]) );
  QDFFS gray_img_reg_9__0__0_ ( .D(n14074), .CK(clk), .Q(gray_img[1152]) );
  QDFFS gray_img_reg_9__2__0_ ( .D(n14065), .CK(clk), .Q(gray_img[1168]) );
  QDFFS gray_img_reg_9__3__0_ ( .D(n14064), .CK(clk), .Q(gray_img[1176]) );
  QDFFS gray_img_reg_9__4__0_ ( .D(n14056), .CK(clk), .Q(gray_img[1184]) );
  QDFFS gray_img_reg_9__5__0_ ( .D(n14055), .CK(clk), .Q(gray_img[1192]) );
  QDFFS gray_img_reg_9__6__0_ ( .D(n14047), .CK(clk), .Q(gray_img[1200]) );
  QDFFS gray_img_reg_9__7__0_ ( .D(n14046), .CK(clk), .Q(gray_img[1208]) );
  QDFFS gray_img_reg_9__8__0_ ( .D(n14038), .CK(clk), .Q(gray_img[1216]) );
  QDFFS gray_img_reg_9__9__0_ ( .D(n14037), .CK(clk), .Q(gray_img[1224]) );
  QDFFS gray_img_reg_9__10__0_ ( .D(n14029), .CK(clk), .Q(gray_img[1232]) );
  QDFFS gray_img_reg_9__11__0_ ( .D(n14028), .CK(clk), .Q(gray_img[1240]) );
  QDFFS gray_img_reg_9__14__0_ ( .D(n14011), .CK(clk), .Q(gray_img[1264]) );
  QDFFS gray_img_reg_9__15__0_ ( .D(n14010), .CK(clk), .Q(gray_img[1272]) );
  QDFFS gray_img_reg_10__1__0_ ( .D(n14001), .CK(clk), .Q(gray_img[1288]) );
  QDFFS gray_img_reg_10__3__0_ ( .D(n13999), .CK(clk), .Q(gray_img[1304]) );
  QDFFS gray_img_reg_10__4__0_ ( .D(n13998), .CK(clk), .Q(gray_img[1312]) );
  QDFFS gray_img_reg_10__6__0_ ( .D(n13996), .CK(clk), .Q(gray_img[1328]) );
  QDFFS gray_img_reg_10__7__0_ ( .D(n13995), .CK(clk), .Q(gray_img[1336]) );
  QDFFS gray_img_reg_10__8__0_ ( .D(n13994), .CK(clk), .Q(gray_img[1344]) );
  QDFFS gray_img_reg_10__10__0_ ( .D(n13992), .CK(clk), .Q(gray_img[1360]) );
  QDFFS gray_img_reg_10__11__0_ ( .D(n13991), .CK(clk), .Q(gray_img[1368]) );
  QDFFS gray_img_reg_10__12__0_ ( .D(n13990), .CK(clk), .Q(gray_img[1376]) );
  QDFFS gray_img_reg_10__13__0_ ( .D(n13989), .CK(clk), .Q(gray_img[1384]) );
  QDFFS gray_img_reg_10__14__0_ ( .D(n13988), .CK(clk), .Q(gray_img[1392]) );
  QDFFS gray_img_reg_10__15__0_ ( .D(n13987), .CK(clk), .Q(gray_img[1400]) );
  QDFFS gray_img_reg_11__0__0_ ( .D(n13986), .CK(clk), .Q(gray_img[1408]) );
  QDFFS gray_img_reg_11__1__0_ ( .D(n13985), .CK(clk), .Q(gray_img[1416]) );
  QDFFS gray_img_reg_11__2__0_ ( .D(n13977), .CK(clk), .Q(gray_img[1424]) );
  QDFFS gray_img_reg_11__3__0_ ( .D(n13976), .CK(clk), .Q(gray_img[1432]) );
  QDFFS gray_img_reg_11__4__0_ ( .D(n13968), .CK(clk), .Q(gray_img[1440]) );
  QDFFS gray_img_reg_11__5__0_ ( .D(n13967), .CK(clk), .Q(gray_img[1448]) );
  QDFFS gray_img_reg_11__6__0_ ( .D(n13959), .CK(clk), .Q(gray_img[1456]) );
  QDFFS gray_img_reg_11__7__0_ ( .D(n13958), .CK(clk), .Q(gray_img[1464]) );
  QDFFS gray_img_reg_11__9__0_ ( .D(n13950), .CK(clk), .Q(gray_img[1480]) );
  QDFFS gray_img_reg_11__10__0_ ( .D(n13943), .CK(clk), .Q(gray_img[1488]) );
  QDFFS gray_img_reg_11__11__0_ ( .D(n13942), .CK(clk), .Q(gray_img[1496]) );
  QDFFS gray_img_reg_11__12__0_ ( .D(n13936), .CK(clk), .Q(gray_img[1504]) );
  QDFFS gray_img_reg_11__13__0_ ( .D(n13935), .CK(clk), .Q(gray_img[1512]) );
  QDFFS gray_img_reg_11__14__0_ ( .D(n13929), .CK(clk), .Q(gray_img[1520]) );
  QDFFS gray_img_reg_11__15__0_ ( .D(n13928), .CK(clk), .Q(gray_img[1528]) );
  QDFFS gray_img_reg_12__0__0_ ( .D(n13923), .CK(clk), .Q(gray_img[1536]) );
  QDFFS gray_img_reg_12__1__0_ ( .D(n13922), .CK(clk), .Q(gray_img[1544]) );
  QDFFS gray_img_reg_12__2__0_ ( .D(n13921), .CK(clk), .Q(gray_img[1552]) );
  QDFFS gray_img_reg_12__3__0_ ( .D(n13920), .CK(clk), .Q(gray_img[1560]) );
  QDFFS gray_img_reg_12__4__0_ ( .D(n13919), .CK(clk), .Q(gray_img[1568]) );
  QDFFS gray_img_reg_12__5__0_ ( .D(n13918), .CK(clk), .Q(gray_img[1576]) );
  QDFFS gray_img_reg_12__6__0_ ( .D(n13917), .CK(clk), .Q(gray_img[1584]) );
  QDFFS gray_img_reg_12__7__0_ ( .D(n13916), .CK(clk), .Q(gray_img[1592]) );
  QDFFS gray_img_reg_12__8__0_ ( .D(n13915), .CK(clk), .Q(gray_img[1600]) );
  QDFFS gray_img_reg_12__9__0_ ( .D(n13914), .CK(clk), .Q(gray_img[1608]) );
  QDFFS gray_img_reg_12__11__0_ ( .D(n13912), .CK(clk), .Q(gray_img[1624]) );
  QDFFS gray_img_reg_12__12__0_ ( .D(n13911), .CK(clk), .Q(gray_img[1632]) );
  QDFFS gray_img_reg_12__13__0_ ( .D(n13910), .CK(clk), .Q(gray_img[1640]) );
  QDFFS gray_img_reg_12__14__0_ ( .D(n13909), .CK(clk), .Q(gray_img[1648]) );
  QDFFS gray_img_reg_13__0__0_ ( .D(n13907), .CK(clk), .Q(gray_img[1664]) );
  QDFFS gray_img_reg_13__1__0_ ( .D(n13906), .CK(clk), .Q(gray_img[1672]) );
  QDFFS gray_img_reg_13__2__0_ ( .D(n13901), .CK(clk), .Q(gray_img[1680]) );
  QDFFS gray_img_reg_13__3__0_ ( .D(n13900), .CK(clk), .Q(gray_img[1688]) );
  QDFFS gray_img_reg_13__4__0_ ( .D(n13895), .CK(clk), .Q(gray_img[1696]) );
  QDFFS gray_img_reg_13__5__0_ ( .D(n13894), .CK(clk), .Q(gray_img[1704]) );
  QDFFS gray_img_reg_13__6__0_ ( .D(n13889), .CK(clk), .Q(gray_img[1712]) );
  QDFFS gray_img_reg_13__7__0_ ( .D(n13888), .CK(clk), .Q(gray_img[1720]) );
  QDFFS gray_img_reg_13__8__0_ ( .D(n13883), .CK(clk), .Q(gray_img[1728]) );
  QDFFS gray_img_reg_13__9__0_ ( .D(n13882), .CK(clk), .Q(gray_img[1736]) );
  QDFFS gray_img_reg_13__10__0_ ( .D(n13877), .CK(clk), .Q(gray_img[1744]) );
  QDFFS gray_img_reg_13__11__0_ ( .D(n13876), .CK(clk), .Q(gray_img[1752]) );
  QDFFS gray_img_reg_13__12__0_ ( .D(n13871), .CK(clk), .Q(gray_img[1760]) );
  QDFFS gray_img_reg_13__13__0_ ( .D(n13870), .CK(clk), .Q(gray_img[1768]) );
  QDFFS gray_img_reg_13__14__0_ ( .D(n13865), .CK(clk), .Q(gray_img[1776]) );
  QDFFS gray_img_reg_13__15__0_ ( .D(n13864), .CK(clk), .Q(gray_img[1784]) );
  QDFFS gray_img_reg_14__0__0_ ( .D(n13859), .CK(clk), .Q(gray_img[1792]) );
  QDFFS gray_img_reg_14__1__0_ ( .D(n13858), .CK(clk), .Q(gray_img[1800]) );
  QDFFS gray_img_reg_14__2__0_ ( .D(n13857), .CK(clk), .Q(gray_img[1808]) );
  QDFFS gray_img_reg_14__4__0_ ( .D(n13855), .CK(clk), .Q(gray_img[1824]) );
  QDFFS gray_img_reg_14__5__0_ ( .D(n13854), .CK(clk), .Q(gray_img[1832]) );
  QDFFS gray_img_reg_14__7__0_ ( .D(n13852), .CK(clk), .Q(gray_img[1848]) );
  QDFFS gray_img_reg_14__8__0_ ( .D(n13851), .CK(clk), .Q(gray_img[1856]) );
  QDFFS gray_img_reg_14__9__0_ ( .D(n13850), .CK(clk), .Q(gray_img[1864]) );
  QDFFS gray_img_reg_14__10__0_ ( .D(n13849), .CK(clk), .Q(gray_img[1872]) );
  QDFFS gray_img_reg_14__11__0_ ( .D(n13848), .CK(clk), .Q(gray_img[1880]) );
  QDFFS gray_img_reg_14__13__0_ ( .D(n13846), .CK(clk), .Q(gray_img[1896]) );
  QDFFS gray_img_reg_15__0__0_ ( .D(n13843), .CK(clk), .Q(gray_img[1920]) );
  QDFFS gray_img_reg_15__1__0_ ( .D(n13842), .CK(clk), .Q(gray_img[1928]) );
  QDFFS gray_img_reg_15__2__0_ ( .D(n13837), .CK(clk), .Q(gray_img[1936]) );
  QDFFS gray_img_reg_15__3__0_ ( .D(n13836), .CK(clk), .Q(gray_img[1944]) );
  QDFFS gray_img_reg_15__5__0_ ( .D(n13831), .CK(clk), .Q(gray_img[1960]) );
  QDFFS gray_img_reg_15__6__0_ ( .D(n13827), .CK(clk), .Q(gray_img[1968]) );
  QDFFS gray_img_reg_15__7__0_ ( .D(n13826), .CK(clk), .Q(gray_img[1976]) );
  QDFFS gray_img_reg_15__9__0_ ( .D(n13822), .CK(clk), .Q(gray_img[1992]) );
  QDFFS gray_img_reg_15__10__0_ ( .D(n13819), .CK(clk), .Q(gray_img[2000]) );
  QDFFS gray_img_reg_15__11__0_ ( .D(n13818), .CK(clk), .Q(gray_img[2008]) );
  QDFFS gray_img_reg_15__12__0_ ( .D(n13816), .CK(clk), .Q(gray_img[2016]) );
  QDFFS gray_img_reg_15__14__0_ ( .D(n13813), .CK(clk), .Q(gray_img[2032]) );
  QDFFS gray_img_reg_15__15__0_ ( .D(n13812), .CK(clk), .Q(gray_img[2040]) );
  QDFFS gray_img_reg_0__4__0_ ( .D(n13810), .CK(clk), .Q(gray_img[32]) );
  QDFFS gray_img_reg_0__6__0_ ( .D(n13808), .CK(clk), .Q(gray_img[48]) );
  QDFFS gray_img_reg_0__7__0_ ( .D(n13807), .CK(clk), .Q(gray_img[56]) );
  QDFFS gray_img_reg_1__4__0_ ( .D(n13804), .CK(clk), .Q(gray_img[160]) );
  QDFFS gray_img_reg_1__5__0_ ( .D(n13803), .CK(clk), .Q(gray_img[168]) );
  QDFFS gray_img_reg_1__6__0_ ( .D(n13794), .CK(clk), .Q(gray_img[176]) );
  QDFFS gray_img_reg_0__3__0_ ( .D(n13792), .CK(clk), .Q(gray_img[24]) );
  QDFFS gray_img_reg_2__4__0_ ( .D(n13782), .CK(clk), .Q(gray_img[288]) );
  QDFFS gray_img_reg_2__7__0_ ( .D(n13779), .CK(clk), .Q(gray_img[312]) );
  QDFFS gray_img_reg_3__4__0_ ( .D(n13774), .CK(clk), .Q(gray_img[416]) );
  QDFFS gray_img_reg_3__5__0_ ( .D(n13773), .CK(clk), .Q(gray_img[424]) );
  QDFFS gray_img_reg_1__2__0_ ( .D(n13772), .CK(clk), .Q(gray_img[144]) );
  QDFFS gray_img_reg_3__6__0_ ( .D(n13764), .CK(clk), .Q(gray_img[432]) );
  QDFFS gray_img_reg_1__3__0_ ( .D(n13762), .CK(clk), .Q(gray_img[152]) );
  QDFFS gray_img_reg_0__1__0_ ( .D(n13754), .CK(clk), .Q(gray_img[8]) );
  QDFFS gray_img_reg_4__1__0_ ( .D(n13745), .CK(clk), .Q(gray_img[520]) );
  QDFFS gray_img_reg_4__2__0_ ( .D(n13744), .CK(clk), .Q(gray_img[528]) );
  QDFFS gray_img_reg_4__3__0_ ( .D(n13743), .CK(clk), .Q(gray_img[536]) );
  QDFFS gray_img_reg_4__4__0_ ( .D(n13742), .CK(clk), .Q(gray_img[544]) );
  QDFFS gray_img_reg_4__6__0_ ( .D(n13740), .CK(clk), .Q(gray_img[560]) );
  QDFFS gray_img_reg_5__0__0_ ( .D(n13738), .CK(clk), .Q(gray_img[640]) );
  QDFFS gray_img_reg_5__1__0_ ( .D(n13737), .CK(clk), .Q(gray_img[648]) );
  QDFFS gray_img_reg_5__3__0_ ( .D(n13727), .CK(clk), .Q(gray_img[664]) );
  QDFFS gray_img_reg_2__1__0_ ( .D(n14267), .CK(clk), .Q(gray_img[264]) );
  QDFFS gray_img_reg_5__4__0_ ( .D(n13726), .CK(clk), .Q(gray_img[672]) );
  QDFFS gray_img_reg_5__5__0_ ( .D(n13725), .CK(clk), .Q(gray_img[680]) );
  QDFFS gray_img_reg_2__2__0_ ( .D(n13784), .CK(clk), .Q(gray_img[272]) );
  QDFFS gray_img_reg_5__6__0_ ( .D(n13724), .CK(clk), .Q(gray_img[688]) );
  QDFFS gray_img_reg_5__7__0_ ( .D(n13723), .CK(clk), .Q(gray_img[696]) );
  QDFFS gray_img_reg_2__3__0_ ( .D(n13783), .CK(clk), .Q(gray_img[280]) );
  QDFFS gray_img_reg_6__0__0_ ( .D(n13722), .CK(clk), .Q(gray_img[768]) );
  QDFFS gray_img_reg_6__1__0_ ( .D(n13721), .CK(clk), .Q(gray_img[776]) );
  QDFFS gray_img_reg_6__2__0_ ( .D(n13720), .CK(clk), .Q(gray_img[784]) );
  QDFFS gray_img_reg_6__3__0_ ( .D(n13719), .CK(clk), .Q(gray_img[792]) );
  QDFFS gray_img_reg_6__4__0_ ( .D(n13718), .CK(clk), .Q(gray_img[800]) );
  QDFFS gray_img_reg_6__6__0_ ( .D(n13716), .CK(clk), .Q(gray_img[816]) );
  QDFFS gray_img_reg_6__7__0_ ( .D(n13715), .CK(clk), .Q(gray_img[824]) );
  QDFFS gray_img_reg_7__0__0_ ( .D(n13714), .CK(clk), .Q(gray_img[896]) );
  QDFFS gray_img_reg_7__1__0_ ( .D(n13713), .CK(clk), .Q(gray_img[904]) );
  QDFFS gray_img_reg_3__0__0_ ( .D(n13778), .CK(clk), .Q(gray_img[384]) );
  QDFFS gray_img_reg_7__2__0_ ( .D(n13712), .CK(clk), .Q(gray_img[912]) );
  QDFFS gray_img_reg_7__3__0_ ( .D(n13711), .CK(clk), .Q(gray_img[920]) );
  QDFFS gray_img_reg_3__1__0_ ( .D(n13777), .CK(clk), .Q(gray_img[392]) );
  QDFFS gray_img_reg_1__0__0_ ( .D(n13806), .CK(clk), .Q(gray_img[128]) );
  QDFFS gray_img_reg_7__4__0_ ( .D(n13710), .CK(clk), .Q(gray_img[928]) );
  QDFFS gray_img_reg_7__5__0_ ( .D(n13709), .CK(clk), .Q(gray_img[936]) );
  QDFFS gray_img_reg_3__2__0_ ( .D(n13776), .CK(clk), .Q(gray_img[400]) );
  QDFFS gray_img_reg_7__6__0_ ( .D(n13708), .CK(clk), .Q(gray_img[944]) );
  QDFFS gray_img_reg_7__7__0_ ( .D(n13707), .CK(clk), .Q(gray_img[952]) );
  QDFFS gray_img_reg_3__3__0_ ( .D(n13775), .CK(clk), .Q(gray_img[408]) );
  QDFFS gray_img_reg_1__1__0_ ( .D(n13805), .CK(clk), .Q(gray_img[136]) );
  QDFFS gray_img_reg_0__0__7_ ( .D(n13613), .CK(clk), .Q(gray_img[7]) );
  QDFFS mem_data_out_reg_shift_0_reg_0__7_ ( .D(n15808), .CK(clk), .Q(
        mem_data_out_reg_shift_0[7]) );
  QDFFS mem_data_out_reg_shift_0_reg_1__7_ ( .D(mem_data_out_reg_shift_0[7]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[15]) );
  QDFFS mem_data_out_reg_shift_0_reg_2__7_ ( .D(mem_data_out_reg_shift_0[15]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[23]) );
  QDFFS mem_data_out_reg_shift_0_reg_3__7_ ( .D(mem_data_out_reg_shift_0[23]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[31]) );
  QDFFS mem_data_out_reg_shift_0_reg_4__7_ ( .D(mem_data_out_reg_shift_0[31]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[39]) );
  QDFFS mem_data_out_reg_shift_0_reg_5__7_ ( .D(mem_data_out_reg_shift_0[39]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[47]) );
  QDFFS mem_data_out_reg_shift_0_reg_6__7_ ( .D(mem_data_out_reg_shift_0[47]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[55]) );
  QDFFS mem_data_out_reg_shift_0_reg_7__7_ ( .D(mem_data_out_reg_shift_0[55]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[63]) );
  QDFFS mem_data_out_reg_shift_0_reg_8__7_ ( .D(mem_data_out_reg_shift_0[63]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[71]) );
  QDFFS mem_data_out_reg_shift_0_reg_9__7_ ( .D(mem_data_out_reg_shift_0[71]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[79]) );
  QDFFS mem_data_out_reg_shift_0_reg_10__7_ ( .D(mem_data_out_reg_shift_0[79]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[87]) );
  QDFFS mem_data_out_reg_shift_0_reg_11__7_ ( .D(mem_data_out_reg_shift_0[87]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[95]) );
  QDFFS mem_data_out_reg_shift_0_reg_12__7_ ( .D(mem_data_out_reg_shift_0[95]), 
        .CK(clk), .Q(mem_data_out_reg_shift_0[103]) );
  QDFFS mem_data_out_reg_shift_0_reg_13__7_ ( .D(mem_data_out_reg_shift_0[103]), .CK(clk), .Q(mem_data_out_reg_shift_0[111]) );
  QDFFS mem_data_out_reg_shift_0_reg_14__7_ ( .D(mem_data_out_reg_shift_0[111]), .CK(clk), .Q(mem_data_out_reg_shift_0[119]) );
  QDFFS mem_data_out_reg_shift_0_reg_15__7_ ( .D(mem_data_out_reg_shift_0[119]), .CK(clk), .Q(mem_data_out_reg_shift_0[127]) );
  QDFFS mem_data_out_reg_shift_1_reg_0__7_ ( .D(n15825), .CK(clk), .Q(
        mem_data_out_reg_shift_1[7]) );
  QDFFS mem_data_out_reg_shift_1_reg_1__7_ ( .D(mem_data_out_reg_shift_1[7]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[15]) );
  QDFFS mem_data_out_reg_shift_1_reg_3__7_ ( .D(mem_data_out_reg_shift_1[23]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[31]) );
  QDFFS mem_data_out_reg_shift_1_reg_4__7_ ( .D(mem_data_out_reg_shift_1[31]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[39]) );
  QDFFS mem_data_out_reg_shift_1_reg_5__7_ ( .D(mem_data_out_reg_shift_1[39]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[47]) );
  QDFFS mem_data_out_reg_shift_1_reg_6__7_ ( .D(mem_data_out_reg_shift_1[47]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[55]) );
  QDFFS mem_data_out_reg_shift_1_reg_7__7_ ( .D(mem_data_out_reg_shift_1[55]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[63]) );
  QDFFS mem_data_out_reg_shift_1_reg_8__7_ ( .D(mem_data_out_reg_shift_1[63]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[71]) );
  QDFFS mem_data_out_reg_shift_1_reg_9__7_ ( .D(mem_data_out_reg_shift_1[71]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[79]) );
  QDFFS mem_data_out_reg_shift_1_reg_10__7_ ( .D(mem_data_out_reg_shift_1[79]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[87]) );
  QDFFS mem_data_out_reg_shift_1_reg_11__7_ ( .D(mem_data_out_reg_shift_1[87]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[95]) );
  QDFFS mem_data_out_reg_shift_1_reg_12__7_ ( .D(mem_data_out_reg_shift_1[95]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[103]) );
  QDFFS mem_data_out_reg_shift_1_reg_13__7_ ( .D(mem_data_out_reg_shift_1[103]), .CK(clk), .Q(mem_data_out_reg_shift_1[111]) );
  QDFFS mem_data_out_reg_shift_1_reg_14__7_ ( .D(mem_data_out_reg_shift_1[111]), .CK(clk), .Q(mem_data_out_reg_shift_1[119]) );
  QDFFS mem_data_out_reg_shift_1_reg_15__7_ ( .D(mem_data_out_reg_shift_1[119]), .CK(clk), .Q(mem_data_out_reg_shift_1[127]) );
  QDFFS mem_data_out_reg_shift_2_reg_0__7_ ( .D(n15833), .CK(clk), .Q(
        mem_data_out_reg_shift_2[7]) );
  QDFFS mem_data_out_reg_shift_2_reg_2__7_ ( .D(mem_data_out_reg_shift_2[15]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[23]) );
  QDFFS mem_data_out_reg_shift_2_reg_3__7_ ( .D(mem_data_out_reg_shift_2[23]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[31]) );
  QDFFS gray_img_reg_15__15__7_ ( .D(n15660), .CK(clk), .Q(gray_img[2047]) );
  QDFFS gray_img_reg_0__8__7_ ( .D(n15659), .CK(clk), .Q(gray_img[71]) );
  QDFFS gray_img_reg_0__9__7_ ( .D(n15658), .CK(clk), .Q(gray_img[79]) );
  QDFFS gray_img_reg_0__10__7_ ( .D(n15657), .CK(clk), .Q(gray_img[87]) );
  QDFFS gray_img_reg_0__11__7_ ( .D(n15656), .CK(clk), .Q(gray_img[95]) );
  QDFFS gray_img_reg_0__12__7_ ( .D(n15655), .CK(clk), .Q(gray_img[103]) );
  QDFFS gray_img_reg_0__13__7_ ( .D(n15654), .CK(clk), .Q(gray_img[111]) );
  QDFFS gray_img_reg_0__14__7_ ( .D(n15653), .CK(clk), .Q(gray_img[119]) );
  QDFFS gray_img_reg_0__15__7_ ( .D(n15652), .CK(clk), .Q(gray_img[127]) );
  QDFFS gray_img_reg_1__8__7_ ( .D(n15651), .CK(clk), .Q(gray_img[199]) );
  QDFFS gray_img_reg_1__9__7_ ( .D(n15650), .CK(clk), .Q(gray_img[207]) );
  QDFFS gray_img_reg_1__10__7_ ( .D(n15649), .CK(clk), .Q(gray_img[215]) );
  QDFFS gray_img_reg_1__11__7_ ( .D(n15648), .CK(clk), .Q(gray_img[223]) );
  QDFFS gray_img_reg_1__12__7_ ( .D(n15647), .CK(clk), .Q(gray_img[231]) );
  QDFFS gray_img_reg_1__13__7_ ( .D(n15646), .CK(clk), .Q(gray_img[239]) );
  QDFFS gray_img_reg_1__14__7_ ( .D(n15645), .CK(clk), .Q(gray_img[247]) );
  QDFFS gray_img_reg_1__15__7_ ( .D(n15644), .CK(clk), .Q(gray_img[255]) );
  QDFFS gray_img_reg_2__8__7_ ( .D(n15643), .CK(clk), .Q(gray_img[327]) );
  QDFFS gray_img_reg_2__9__7_ ( .D(n15642), .CK(clk), .Q(gray_img[335]) );
  QDFFS gray_img_reg_2__10__7_ ( .D(n15641), .CK(clk), .Q(gray_img[343]) );
  QDFFS gray_img_reg_2__11__7_ ( .D(n15640), .CK(clk), .Q(gray_img[351]) );
  QDFFS gray_img_reg_2__12__7_ ( .D(n15639), .CK(clk), .Q(gray_img[359]) );
  QDFFS gray_img_reg_2__13__7_ ( .D(n15638), .CK(clk), .Q(gray_img[367]) );
  QDFFS gray_img_reg_2__14__7_ ( .D(n15637), .CK(clk), .Q(gray_img[375]) );
  QDFFS gray_img_reg_2__15__7_ ( .D(n15636), .CK(clk), .Q(gray_img[383]) );
  QDFFS gray_img_reg_3__8__7_ ( .D(n15635), .CK(clk), .Q(gray_img[455]) );
  QDFFS gray_img_reg_3__9__7_ ( .D(n15634), .CK(clk), .Q(gray_img[463]) );
  QDFFS gray_img_reg_3__10__7_ ( .D(n15633), .CK(clk), .Q(gray_img[471]) );
  QDFFS gray_img_reg_3__11__7_ ( .D(n15632), .CK(clk), .Q(gray_img[479]) );
  QDFFS gray_img_reg_3__12__7_ ( .D(n15631), .CK(clk), .Q(gray_img[487]) );
  QDFFS gray_img_reg_3__13__7_ ( .D(n15630), .CK(clk), .Q(gray_img[495]) );
  QDFFS gray_img_reg_3__14__7_ ( .D(n15629), .CK(clk), .Q(gray_img[503]) );
  QDFFS gray_img_reg_3__15__7_ ( .D(n15628), .CK(clk), .Q(gray_img[511]) );
  QDFFS gray_img_reg_4__8__7_ ( .D(n15627), .CK(clk), .Q(gray_img[583]) );
  QDFFS gray_img_reg_4__9__7_ ( .D(n15626), .CK(clk), .Q(gray_img[591]) );
  QDFFS gray_img_reg_4__10__7_ ( .D(n15625), .CK(clk), .Q(gray_img[599]) );
  QDFFS gray_img_reg_4__11__7_ ( .D(n15624), .CK(clk), .Q(gray_img[607]) );
  QDFFS gray_img_reg_4__12__7_ ( .D(n15623), .CK(clk), .Q(gray_img[615]) );
  QDFFS gray_img_reg_4__13__7_ ( .D(n15622), .CK(clk), .Q(gray_img[623]) );
  QDFFS gray_img_reg_4__14__7_ ( .D(n15621), .CK(clk), .Q(gray_img[631]) );
  QDFFS gray_img_reg_4__15__7_ ( .D(n15620), .CK(clk), .Q(gray_img[639]) );
  QDFFS gray_img_reg_5__8__7_ ( .D(n15619), .CK(clk), .Q(gray_img[711]) );
  QDFFS gray_img_reg_5__9__7_ ( .D(n15618), .CK(clk), .Q(gray_img[719]) );
  QDFFS gray_img_reg_5__10__7_ ( .D(n15617), .CK(clk), .Q(gray_img[727]) );
  QDFFS gray_img_reg_5__11__7_ ( .D(n15616), .CK(clk), .Q(gray_img[735]) );
  QDFFS gray_img_reg_5__12__7_ ( .D(n15615), .CK(clk), .Q(gray_img[743]) );
  QDFFS gray_img_reg_5__13__7_ ( .D(n15614), .CK(clk), .Q(gray_img[751]) );
  QDFFS gray_img_reg_5__14__7_ ( .D(n15613), .CK(clk), .Q(gray_img[759]) );
  QDFFS gray_img_reg_5__15__7_ ( .D(n15612), .CK(clk), .Q(gray_img[767]) );
  QDFFS gray_img_reg_6__8__7_ ( .D(n15611), .CK(clk), .Q(gray_img[839]) );
  QDFFS gray_img_reg_6__9__7_ ( .D(n15610), .CK(clk), .Q(gray_img[847]) );
  QDFFS gray_img_reg_6__10__7_ ( .D(n15609), .CK(clk), .Q(gray_img[855]) );
  QDFFS gray_img_reg_6__11__7_ ( .D(n15608), .CK(clk), .Q(gray_img[863]) );
  QDFFS gray_img_reg_6__12__7_ ( .D(n15607), .CK(clk), .Q(gray_img[871]) );
  QDFFS gray_img_reg_6__13__7_ ( .D(n15606), .CK(clk), .Q(gray_img[879]) );
  QDFFS gray_img_reg_6__14__7_ ( .D(n15605), .CK(clk), .Q(gray_img[887]) );
  QDFFS gray_img_reg_6__15__7_ ( .D(n15604), .CK(clk), .Q(gray_img[895]) );
  QDFFS gray_img_reg_7__8__7_ ( .D(n15603), .CK(clk), .Q(gray_img[967]) );
  QDFFS gray_img_reg_7__9__7_ ( .D(n15602), .CK(clk), .Q(gray_img[975]) );
  QDFFS gray_img_reg_7__10__7_ ( .D(n15601), .CK(clk), .Q(gray_img[983]) );
  QDFFS gray_img_reg_7__11__7_ ( .D(n15600), .CK(clk), .Q(gray_img[991]) );
  QDFFS gray_img_reg_7__12__7_ ( .D(n15599), .CK(clk), .Q(gray_img[999]) );
  QDFFS gray_img_reg_7__13__7_ ( .D(n15598), .CK(clk), .Q(gray_img[1007]) );
  QDFFS gray_img_reg_7__14__7_ ( .D(n15597), .CK(clk), .Q(gray_img[1015]) );
  QDFFS gray_img_reg_7__15__7_ ( .D(n15596), .CK(clk), .Q(gray_img[1023]) );
  QDFFS gray_img_reg_8__0__7_ ( .D(n15595), .CK(clk), .Q(gray_img[1031]) );
  QDFFS gray_img_reg_8__1__7_ ( .D(n15594), .CK(clk), .Q(gray_img[1039]) );
  QDFFS gray_img_reg_8__2__7_ ( .D(n15593), .CK(clk), .Q(gray_img[1047]) );
  QDFFS gray_img_reg_8__3__7_ ( .D(n15592), .CK(clk), .Q(gray_img[1055]) );
  QDFFS gray_img_reg_8__4__7_ ( .D(n15591), .CK(clk), .Q(gray_img[1063]) );
  QDFFS gray_img_reg_8__5__7_ ( .D(n15590), .CK(clk), .Q(gray_img[1071]) );
  QDFFS gray_img_reg_8__6__7_ ( .D(n15589), .CK(clk), .Q(gray_img[1079]) );
  QDFFS gray_img_reg_8__7__7_ ( .D(n15588), .CK(clk), .Q(gray_img[1087]) );
  QDFFS gray_img_reg_8__8__7_ ( .D(n15587), .CK(clk), .Q(gray_img[1095]) );
  QDFFS gray_img_reg_8__9__7_ ( .D(n15586), .CK(clk), .Q(gray_img[1103]) );
  QDFFS gray_img_reg_8__10__7_ ( .D(n15585), .CK(clk), .Q(gray_img[1111]) );
  QDFFS gray_img_reg_8__11__7_ ( .D(n15584), .CK(clk), .Q(gray_img[1119]) );
  QDFFS gray_img_reg_8__12__7_ ( .D(n15583), .CK(clk), .Q(gray_img[1127]) );
  QDFFS gray_img_reg_8__13__7_ ( .D(n15582), .CK(clk), .Q(gray_img[1135]) );
  QDFFS gray_img_reg_8__14__7_ ( .D(n15581), .CK(clk), .Q(gray_img[1143]) );
  QDFFS gray_img_reg_8__15__7_ ( .D(n15580), .CK(clk), .Q(gray_img[1151]) );
  QDFFS gray_img_reg_9__0__7_ ( .D(n15579), .CK(clk), .Q(gray_img[1159]) );
  QDFFS gray_img_reg_9__1__7_ ( .D(n15578), .CK(clk), .Q(gray_img[1167]) );
  QDFFS gray_img_reg_9__2__7_ ( .D(n15577), .CK(clk), .Q(gray_img[1175]) );
  QDFFS gray_img_reg_9__3__7_ ( .D(n15576), .CK(clk), .Q(gray_img[1183]) );
  QDFFS gray_img_reg_9__4__7_ ( .D(n15575), .CK(clk), .Q(gray_img[1191]) );
  QDFFS gray_img_reg_9__5__7_ ( .D(n15574), .CK(clk), .Q(gray_img[1199]) );
  QDFFS gray_img_reg_9__6__7_ ( .D(n15573), .CK(clk), .Q(gray_img[1207]) );
  QDFFS gray_img_reg_9__7__7_ ( .D(n15572), .CK(clk), .Q(gray_img[1215]) );
  QDFFS gray_img_reg_9__8__7_ ( .D(n15571), .CK(clk), .Q(gray_img[1223]) );
  QDFFS gray_img_reg_9__9__7_ ( .D(n15570), .CK(clk), .Q(gray_img[1231]) );
  QDFFS gray_img_reg_9__10__7_ ( .D(n15569), .CK(clk), .Q(gray_img[1239]) );
  QDFFS gray_img_reg_9__11__7_ ( .D(n15568), .CK(clk), .Q(gray_img[1247]) );
  QDFFS gray_img_reg_9__12__7_ ( .D(n15567), .CK(clk), .Q(gray_img[1255]) );
  QDFFS gray_img_reg_9__13__7_ ( .D(n15566), .CK(clk), .Q(gray_img[1263]) );
  QDFFS gray_img_reg_9__14__7_ ( .D(n15565), .CK(clk), .Q(gray_img[1271]) );
  QDFFS gray_img_reg_9__15__7_ ( .D(n15564), .CK(clk), .Q(gray_img[1279]) );
  QDFFS gray_img_reg_10__0__7_ ( .D(n15563), .CK(clk), .Q(gray_img[1287]) );
  QDFFS gray_img_reg_10__1__7_ ( .D(n15562), .CK(clk), .Q(gray_img[1295]) );
  QDFFS gray_img_reg_10__2__7_ ( .D(n15561), .CK(clk), .Q(gray_img[1303]) );
  QDFFS gray_img_reg_10__3__7_ ( .D(n15560), .CK(clk), .Q(gray_img[1311]) );
  QDFFS gray_img_reg_10__4__7_ ( .D(n15559), .CK(clk), .Q(gray_img[1319]) );
  QDFFS gray_img_reg_10__5__7_ ( .D(n15558), .CK(clk), .Q(gray_img[1327]) );
  QDFFS gray_img_reg_10__6__7_ ( .D(n15557), .CK(clk), .Q(gray_img[1335]) );
  QDFFS gray_img_reg_10__7__7_ ( .D(n15556), .CK(clk), .Q(gray_img[1343]) );
  QDFFS gray_img_reg_10__8__7_ ( .D(n15555), .CK(clk), .Q(gray_img[1351]) );
  QDFFS gray_img_reg_10__9__7_ ( .D(n15554), .CK(clk), .Q(gray_img[1359]) );
  QDFFS gray_img_reg_10__10__7_ ( .D(n15553), .CK(clk), .Q(gray_img[1367]) );
  QDFFS gray_img_reg_10__11__7_ ( .D(n15552), .CK(clk), .Q(gray_img[1375]) );
  QDFFS gray_img_reg_10__12__7_ ( .D(n15551), .CK(clk), .Q(gray_img[1383]) );
  QDFFS gray_img_reg_10__13__7_ ( .D(n15550), .CK(clk), .Q(gray_img[1391]) );
  QDFFS gray_img_reg_10__14__7_ ( .D(n15549), .CK(clk), .Q(gray_img[1399]) );
  QDFFS gray_img_reg_10__15__7_ ( .D(n15548), .CK(clk), .Q(gray_img[1407]) );
  QDFFS gray_img_reg_11__0__7_ ( .D(n15547), .CK(clk), .Q(gray_img[1415]) );
  QDFFS gray_img_reg_11__1__7_ ( .D(n15546), .CK(clk), .Q(gray_img[1423]) );
  QDFFS gray_img_reg_11__2__7_ ( .D(n15545), .CK(clk), .Q(gray_img[1431]) );
  QDFFS gray_img_reg_11__3__7_ ( .D(n15544), .CK(clk), .Q(gray_img[1439]) );
  QDFFS gray_img_reg_11__4__7_ ( .D(n15543), .CK(clk), .Q(gray_img[1447]) );
  QDFFS gray_img_reg_11__5__7_ ( .D(n15542), .CK(clk), .Q(gray_img[1455]) );
  QDFFS gray_img_reg_11__6__7_ ( .D(n15541), .CK(clk), .Q(gray_img[1463]) );
  QDFFS gray_img_reg_11__7__7_ ( .D(n15540), .CK(clk), .Q(gray_img[1471]) );
  QDFFS gray_img_reg_11__8__7_ ( .D(n15539), .CK(clk), .Q(gray_img[1479]) );
  QDFFS gray_img_reg_11__9__7_ ( .D(n15538), .CK(clk), .Q(gray_img[1487]) );
  QDFFS gray_img_reg_11__10__7_ ( .D(n15537), .CK(clk), .Q(gray_img[1495]) );
  QDFFS gray_img_reg_11__11__7_ ( .D(n15536), .CK(clk), .Q(gray_img[1503]) );
  QDFFS gray_img_reg_11__12__7_ ( .D(n15535), .CK(clk), .Q(gray_img[1511]) );
  QDFFS gray_img_reg_11__13__7_ ( .D(n15534), .CK(clk), .Q(gray_img[1519]) );
  QDFFS gray_img_reg_11__14__7_ ( .D(n15533), .CK(clk), .Q(gray_img[1527]) );
  QDFFS gray_img_reg_11__15__7_ ( .D(n15532), .CK(clk), .Q(gray_img[1535]) );
  QDFFS gray_img_reg_12__0__7_ ( .D(n15531), .CK(clk), .Q(gray_img[1543]) );
  QDFFS gray_img_reg_12__1__7_ ( .D(n15530), .CK(clk), .Q(gray_img[1551]) );
  QDFFS gray_img_reg_12__2__7_ ( .D(n15529), .CK(clk), .Q(gray_img[1559]) );
  QDFFS gray_img_reg_12__3__7_ ( .D(n15528), .CK(clk), .Q(gray_img[1567]) );
  QDFFS gray_img_reg_12__4__7_ ( .D(n15527), .CK(clk), .Q(gray_img[1575]) );
  QDFFS gray_img_reg_12__5__7_ ( .D(n15526), .CK(clk), .Q(gray_img[1583]) );
  QDFFS gray_img_reg_12__6__7_ ( .D(n15525), .CK(clk), .Q(gray_img[1591]) );
  QDFFS gray_img_reg_12__7__7_ ( .D(n15524), .CK(clk), .Q(gray_img[1599]) );
  QDFFS gray_img_reg_12__8__7_ ( .D(n15523), .CK(clk), .Q(gray_img[1607]) );
  QDFFS gray_img_reg_12__9__7_ ( .D(n15522), .CK(clk), .Q(gray_img[1615]) );
  QDFFS gray_img_reg_12__10__7_ ( .D(n15521), .CK(clk), .Q(gray_img[1623]) );
  QDFFS gray_img_reg_12__11__7_ ( .D(n15520), .CK(clk), .Q(gray_img[1631]) );
  QDFFS gray_img_reg_12__12__7_ ( .D(n15519), .CK(clk), .Q(gray_img[1639]) );
  QDFFS gray_img_reg_12__13__7_ ( .D(n15518), .CK(clk), .Q(gray_img[1647]) );
  QDFFS gray_img_reg_12__14__7_ ( .D(n15517), .CK(clk), .Q(gray_img[1655]) );
  QDFFS gray_img_reg_12__15__7_ ( .D(n15516), .CK(clk), .Q(gray_img[1663]) );
  QDFFS gray_img_reg_13__0__7_ ( .D(n15515), .CK(clk), .Q(gray_img[1671]) );
  QDFFS gray_img_reg_13__1__7_ ( .D(n15514), .CK(clk), .Q(gray_img[1679]) );
  QDFFS gray_img_reg_13__2__7_ ( .D(n15513), .CK(clk), .Q(gray_img[1687]) );
  QDFFS gray_img_reg_13__3__7_ ( .D(n15512), .CK(clk), .Q(gray_img[1695]) );
  QDFFS gray_img_reg_13__4__7_ ( .D(n15511), .CK(clk), .Q(gray_img[1703]) );
  QDFFS gray_img_reg_13__5__7_ ( .D(n15510), .CK(clk), .Q(gray_img[1711]) );
  QDFFS gray_img_reg_13__6__7_ ( .D(n15509), .CK(clk), .Q(gray_img[1719]) );
  QDFFS gray_img_reg_13__7__7_ ( .D(n15508), .CK(clk), .Q(gray_img[1727]) );
  QDFFS gray_img_reg_13__8__7_ ( .D(n15507), .CK(clk), .Q(gray_img[1735]) );
  QDFFS gray_img_reg_13__9__7_ ( .D(n15506), .CK(clk), .Q(gray_img[1743]) );
  QDFFS gray_img_reg_13__10__7_ ( .D(n15505), .CK(clk), .Q(gray_img[1751]) );
  QDFFS gray_img_reg_13__11__7_ ( .D(n15504), .CK(clk), .Q(gray_img[1759]) );
  QDFFS gray_img_reg_13__12__7_ ( .D(n15503), .CK(clk), .Q(gray_img[1767]) );
  QDFFS gray_img_reg_13__13__7_ ( .D(n15502), .CK(clk), .Q(gray_img[1775]) );
  QDFFS gray_img_reg_13__14__7_ ( .D(n15501), .CK(clk), .Q(gray_img[1783]) );
  QDFFS gray_img_reg_13__15__7_ ( .D(n15500), .CK(clk), .Q(gray_img[1791]) );
  QDFFS gray_img_reg_14__0__7_ ( .D(n15499), .CK(clk), .Q(gray_img[1799]) );
  QDFFS gray_img_reg_14__1__7_ ( .D(n15498), .CK(clk), .Q(gray_img[1807]) );
  QDFFS gray_img_reg_14__2__7_ ( .D(n15497), .CK(clk), .Q(gray_img[1815]) );
  QDFFS gray_img_reg_14__3__7_ ( .D(n15496), .CK(clk), .Q(gray_img[1823]) );
  QDFFS gray_img_reg_14__4__7_ ( .D(n15495), .CK(clk), .Q(gray_img[1831]) );
  QDFFS gray_img_reg_14__5__7_ ( .D(n15494), .CK(clk), .Q(gray_img[1839]) );
  QDFFS gray_img_reg_14__6__7_ ( .D(n15493), .CK(clk), .Q(gray_img[1847]) );
  QDFFS gray_img_reg_14__7__7_ ( .D(n15492), .CK(clk), .Q(gray_img[1855]) );
  QDFFS gray_img_reg_14__8__7_ ( .D(n15491), .CK(clk), .Q(gray_img[1863]) );
  QDFFS gray_img_reg_14__9__7_ ( .D(n15490), .CK(clk), .Q(gray_img[1871]) );
  QDFFS gray_img_reg_14__10__7_ ( .D(n15489), .CK(clk), .Q(gray_img[1879]) );
  QDFFS gray_img_reg_14__11__7_ ( .D(n15488), .CK(clk), .Q(gray_img[1887]) );
  QDFFS gray_img_reg_14__12__7_ ( .D(n15487), .CK(clk), .Q(gray_img[1895]) );
  QDFFS gray_img_reg_14__13__7_ ( .D(n15486), .CK(clk), .Q(gray_img[1903]) );
  QDFFS gray_img_reg_14__14__7_ ( .D(n15485), .CK(clk), .Q(gray_img[1911]) );
  QDFFS gray_img_reg_14__15__7_ ( .D(n15484), .CK(clk), .Q(gray_img[1919]) );
  QDFFS gray_img_reg_15__0__7_ ( .D(n15483), .CK(clk), .Q(gray_img[1927]) );
  QDFFS gray_img_reg_15__1__7_ ( .D(n15482), .CK(clk), .Q(gray_img[1935]) );
  QDFFS gray_img_reg_15__2__7_ ( .D(n15481), .CK(clk), .Q(gray_img[1943]) );
  QDFFS gray_img_reg_15__3__7_ ( .D(n15480), .CK(clk), .Q(gray_img[1951]) );
  QDFFS gray_img_reg_15__4__7_ ( .D(n15479), .CK(clk), .Q(gray_img[1959]) );
  QDFFS gray_img_reg_15__5__7_ ( .D(n15478), .CK(clk), .Q(gray_img[1967]) );
  QDFFS gray_img_reg_15__6__7_ ( .D(n15477), .CK(clk), .Q(gray_img[1975]) );
  QDFFS gray_img_reg_15__7__7_ ( .D(n15476), .CK(clk), .Q(gray_img[1983]) );
  QDFFS gray_img_reg_15__8__7_ ( .D(n15475), .CK(clk), .Q(gray_img[1991]) );
  QDFFS gray_img_reg_15__9__7_ ( .D(n15474), .CK(clk), .Q(gray_img[1999]) );
  QDFFS gray_img_reg_15__10__7_ ( .D(n15473), .CK(clk), .Q(gray_img[2007]) );
  QDFFS gray_img_reg_15__11__7_ ( .D(n15472), .CK(clk), .Q(gray_img[2015]) );
  QDFFS gray_img_reg_15__12__7_ ( .D(n15471), .CK(clk), .Q(gray_img[2023]) );
  QDFFS gray_img_reg_15__13__7_ ( .D(n15470), .CK(clk), .Q(gray_img[2031]) );
  QDFFS gray_img_reg_15__14__7_ ( .D(n15469), .CK(clk), .Q(gray_img[2039]) );
  QDFFS gray_img_reg_7__7__7_ ( .D(n15468), .CK(clk), .Q(gray_img[959]) );
  QDFFS gray_img_reg_0__4__7_ ( .D(n14250), .CK(clk), .Q(gray_img[39]) );
  QDFFS gray_img_reg_0__5__7_ ( .D(n14241), .CK(clk), .Q(gray_img[47]) );
  QDFFS gray_img_reg_0__6__7_ ( .D(n14232), .CK(clk), .Q(gray_img[55]) );
  QDFFS gray_img_reg_0__7__7_ ( .D(n14223), .CK(clk), .Q(gray_img[63]) );
  QDFFS gray_img_reg_1__4__7_ ( .D(n14206), .CK(clk), .Q(gray_img[167]) );
  QDFFS gray_img_reg_1__5__7_ ( .D(n14197), .CK(clk), .Q(gray_img[175]) );
  QDFFS gray_img_reg_1__6__7_ ( .D(n14188), .CK(clk), .Q(gray_img[183]) );
  QDFFS gray_img_reg_1__7__7_ ( .D(n14179), .CK(clk), .Q(gray_img[191]) );
  QDFFS gray_img_reg_2__4__7_ ( .D(n14162), .CK(clk), .Q(gray_img[295]) );
  QDFFS gray_img_reg_2__5__7_ ( .D(n14153), .CK(clk), .Q(gray_img[303]) );
  QDFFS gray_img_reg_2__6__7_ ( .D(n14144), .CK(clk), .Q(gray_img[311]) );
  QDFFS gray_img_reg_2__7__7_ ( .D(n14135), .CK(clk), .Q(gray_img[319]) );
  QDFFS gray_img_reg_3__4__7_ ( .D(n14118), .CK(clk), .Q(gray_img[423]) );
  QDFFS gray_img_reg_3__5__7_ ( .D(n14109), .CK(clk), .Q(gray_img[431]) );
  QDFFS gray_img_reg_3__6__7_ ( .D(n14100), .CK(clk), .Q(gray_img[439]) );
  QDFFS gray_img_reg_3__7__7_ ( .D(n14091), .CK(clk), .Q(gray_img[447]) );
  QDFFS gray_img_reg_4__0__7_ ( .D(n14066), .CK(clk), .Q(gray_img[519]) );
  QDFFS gray_img_reg_4__1__7_ ( .D(n14057), .CK(clk), .Q(gray_img[527]) );
  QDFFS gray_img_reg_4__2__7_ ( .D(n14048), .CK(clk), .Q(gray_img[535]) );
  QDFFS gray_img_reg_4__3__7_ ( .D(n14039), .CK(clk), .Q(gray_img[543]) );
  QDFFS gray_img_reg_4__4__7_ ( .D(n14030), .CK(clk), .Q(gray_img[551]) );
  QDFFS gray_img_reg_4__5__7_ ( .D(n14021), .CK(clk), .Q(gray_img[559]) );
  QDFFS gray_img_reg_4__6__7_ ( .D(n14012), .CK(clk), .Q(gray_img[567]) );
  QDFFS gray_img_reg_4__7__7_ ( .D(n14003), .CK(clk), .Q(gray_img[575]) );
  QDFFS gray_img_reg_5__0__7_ ( .D(n13978), .CK(clk), .Q(gray_img[647]) );
  QDFFS gray_img_reg_5__1__7_ ( .D(n13969), .CK(clk), .Q(gray_img[655]) );
  QDFFS gray_img_reg_5__2__7_ ( .D(n13960), .CK(clk), .Q(gray_img[663]) );
  QDFFS gray_img_reg_5__3__7_ ( .D(n13952), .CK(clk), .Q(gray_img[671]) );
  QDFFS gray_img_reg_5__4__7_ ( .D(n13944), .CK(clk), .Q(gray_img[679]) );
  QDFFS gray_img_reg_5__5__7_ ( .D(n13937), .CK(clk), .Q(gray_img[687]) );
  QDFFS gray_img_reg_5__6__7_ ( .D(n13930), .CK(clk), .Q(gray_img[695]) );
  QDFFS gray_img_reg_5__7__7_ ( .D(n13924), .CK(clk), .Q(gray_img[703]) );
  QDFFS gray_img_reg_6__0__7_ ( .D(n13902), .CK(clk), .Q(gray_img[775]) );
  QDFFS gray_img_reg_6__1__7_ ( .D(n13896), .CK(clk), .Q(gray_img[783]) );
  QDFFS gray_img_reg_6__2__7_ ( .D(n13890), .CK(clk), .Q(gray_img[791]) );
  QDFFS gray_img_reg_6__3__7_ ( .D(n13884), .CK(clk), .Q(gray_img[799]) );
  QDFFS gray_img_reg_6__4__7_ ( .D(n13878), .CK(clk), .Q(gray_img[807]) );
  QDFFS gray_img_reg_6__5__7_ ( .D(n13872), .CK(clk), .Q(gray_img[815]) );
  QDFFS gray_img_reg_6__6__7_ ( .D(n13866), .CK(clk), .Q(gray_img[823]) );
  QDFFS gray_img_reg_6__7__7_ ( .D(n13860), .CK(clk), .Q(gray_img[831]) );
  QDFFS gray_img_reg_7__0__7_ ( .D(n13838), .CK(clk), .Q(gray_img[903]) );
  QDFFS gray_img_reg_7__1__7_ ( .D(n13833), .CK(clk), .Q(gray_img[911]) );
  QDFFS gray_img_reg_7__2__7_ ( .D(n13828), .CK(clk), .Q(gray_img[919]) );
  QDFFS gray_img_reg_7__3__7_ ( .D(n13824), .CK(clk), .Q(gray_img[927]) );
  QDFFS gray_img_reg_3__1__7_ ( .D(n15070), .CK(clk), .Q(gray_img[399]) );
  QDFFS gray_img_reg_7__4__7_ ( .D(n13820), .CK(clk), .Q(gray_img[935]) );
  QDFFS gray_img_reg_7__5__7_ ( .D(n13817), .CK(clk), .Q(gray_img[943]) );
  QDFFS gray_img_reg_7__6__7_ ( .D(n13814), .CK(clk), .Q(gray_img[951]) );
  QDFFS gray_img_reg_3__3__7_ ( .D(n15467), .CK(clk), .Q(gray_img[415]) );
  QDFFS gray_img_reg_0__2__7_ ( .D(n13795), .CK(clk), .Q(gray_img[23]) );
  QDFFS gray_img_reg_0__3__7_ ( .D(n13785), .CK(clk), .Q(gray_img[31]) );
  QDFFS gray_img_reg_1__2__7_ ( .D(n13765), .CK(clk), .Q(gray_img[151]) );
  QDFFS gray_img_reg_1__3__7_ ( .D(n13755), .CK(clk), .Q(gray_img[159]) );
  QDFFS gray_img_reg_0__1__7_ ( .D(n13747), .CK(clk), .Q(gray_img[15]) );
  QDFFS gray_img_reg_2__0__7_ ( .D(n13729), .CK(clk), .Q(gray_img[263]) );
  QDFFS gray_img_reg_2__1__7_ ( .D(n13700), .CK(clk), .Q(gray_img[271]) );
  QDFFS gray_img_reg_2__2__7_ ( .D(n13674), .CK(clk), .Q(gray_img[279]) );
  QDFFS gray_img_reg_2__3__7_ ( .D(n13651), .CK(clk), .Q(gray_img[287]) );
  QDFFS gray_img_reg_3__0__7_ ( .D(n13631), .CK(clk), .Q(gray_img[391]) );
  QDFFS gray_img_reg_1__0__7_ ( .D(n13622), .CK(clk), .Q(gray_img[135]) );
  QDFFS gray_img_reg_3__2__7_ ( .D(n13616), .CK(clk), .Q(gray_img[407]) );
  QDFFS gray_img_reg_1__1__7_ ( .D(n15466), .CK(clk), .Q(gray_img[143]) );
  QDFFS template_reg_reg_0__0__0_ ( .D(n15732), .CK(clk), .Q(template_reg[0])
         );
  QDFFS template_reg_reg_0__0__1_ ( .D(n15731), .CK(clk), .Q(template_reg[1])
         );
  QDFFS template_reg_reg_0__0__2_ ( .D(n15730), .CK(clk), .Q(template_reg[2])
         );
  QDFFS template_reg_reg_0__0__3_ ( .D(n15729), .CK(clk), .Q(template_reg[3])
         );
  QDFFS template_reg_reg_0__0__4_ ( .D(n15728), .CK(clk), .Q(template_reg[4])
         );
  QDFFS template_reg_reg_0__0__5_ ( .D(n15727), .CK(clk), .Q(template_reg[5])
         );
  QDFFS template_reg_reg_0__0__6_ ( .D(n15726), .CK(clk), .Q(template_reg[6])
         );
  QDFFS template_reg_reg_0__0__7_ ( .D(n15725), .CK(clk), .Q(template_reg[7])
         );
  QDFFS template_reg_reg_0__1__0_ ( .D(n15724), .CK(clk), .Q(template_reg[8])
         );
  QDFFS template_reg_reg_0__1__1_ ( .D(n15723), .CK(clk), .Q(template_reg[9])
         );
  QDFFS template_reg_reg_0__1__2_ ( .D(n15722), .CK(clk), .Q(template_reg[10])
         );
  QDFFS template_reg_reg_0__1__3_ ( .D(n15721), .CK(clk), .Q(template_reg[11])
         );
  QDFFS template_reg_reg_0__1__4_ ( .D(n15720), .CK(clk), .Q(template_reg[12])
         );
  QDFFS template_reg_reg_0__1__5_ ( .D(n15719), .CK(clk), .Q(template_reg[13])
         );
  QDFFS template_reg_reg_0__1__6_ ( .D(n15718), .CK(clk), .Q(template_reg[14])
         );
  QDFFS template_reg_reg_0__1__7_ ( .D(n15717), .CK(clk), .Q(template_reg[15])
         );
  QDFFS template_reg_reg_0__2__0_ ( .D(n15716), .CK(clk), .Q(template_reg[16])
         );
  QDFFS template_reg_reg_0__2__1_ ( .D(n15715), .CK(clk), .Q(template_reg[17])
         );
  QDFFS template_reg_reg_0__2__2_ ( .D(n15714), .CK(clk), .Q(template_reg[18])
         );
  QDFFS template_reg_reg_0__2__3_ ( .D(n15713), .CK(clk), .Q(template_reg[19])
         );
  QDFFS template_reg_reg_0__2__4_ ( .D(n15712), .CK(clk), .Q(template_reg[20])
         );
  QDFFS template_reg_reg_0__2__5_ ( .D(n15711), .CK(clk), .Q(template_reg[21])
         );
  QDFFS template_reg_reg_0__2__6_ ( .D(n15710), .CK(clk), .Q(template_reg[22])
         );
  QDFFS template_reg_reg_0__2__7_ ( .D(n15709), .CK(clk), .Q(template_reg[23])
         );
  QDFFS template_reg_reg_2__0__0_ ( .D(n15684), .CK(clk), .Q(template_reg[48])
         );
  QDFFS template_reg_reg_2__0__1_ ( .D(n15683), .CK(clk), .Q(template_reg[49])
         );
  QDFFS template_reg_reg_2__0__2_ ( .D(n15682), .CK(clk), .Q(template_reg[50])
         );
  QDFFS template_reg_reg_2__0__3_ ( .D(n15681), .CK(clk), .Q(template_reg[51])
         );
  QDFFS template_reg_reg_2__0__4_ ( .D(n15680), .CK(clk), .Q(template_reg[52])
         );
  QDFFS template_reg_reg_2__0__5_ ( .D(n15679), .CK(clk), .Q(template_reg[53])
         );
  QDFFS template_reg_reg_2__0__6_ ( .D(n15678), .CK(clk), .Q(template_reg[54])
         );
  QDFFS template_reg_reg_2__0__7_ ( .D(n15677), .CK(clk), .Q(template_reg[55])
         );
  QDFFS template_reg_reg_2__1__0_ ( .D(n15676), .CK(clk), .Q(template_reg[56])
         );
  QDFFS template_reg_reg_2__1__1_ ( .D(n15675), .CK(clk), .Q(template_reg[57])
         );
  QDFFS template_reg_reg_2__1__2_ ( .D(n15674), .CK(clk), .Q(template_reg[58])
         );
  QDFFS template_reg_reg_2__1__3_ ( .D(n15673), .CK(clk), .Q(template_reg[59])
         );
  QDFFS template_reg_reg_2__1__4_ ( .D(n15672), .CK(clk), .Q(template_reg[60])
         );
  QDFFS template_reg_reg_2__1__5_ ( .D(n15671), .CK(clk), .Q(template_reg[61])
         );
  QDFFS template_reg_reg_2__1__6_ ( .D(n15670), .CK(clk), .Q(template_reg[62])
         );
  QDFFS template_reg_reg_2__1__7_ ( .D(n15669), .CK(clk), .Q(template_reg[63])
         );
  QDFFS template_reg_reg_2__2__0_ ( .D(n15668), .CK(clk), .Q(template_reg[64])
         );
  QDFFS template_reg_reg_2__2__1_ ( .D(n15667), .CK(clk), .Q(template_reg[65])
         );
  QDFFS template_reg_reg_2__2__2_ ( .D(n15666), .CK(clk), .Q(template_reg[66])
         );
  QDFFS template_reg_reg_2__2__3_ ( .D(n15665), .CK(clk), .Q(template_reg[67])
         );
  QDFFS template_reg_reg_2__2__4_ ( .D(n15664), .CK(clk), .Q(template_reg[68])
         );
  QDFFS template_reg_reg_2__2__5_ ( .D(n15663), .CK(clk), .Q(template_reg[69])
         );
  QDFFS template_reg_reg_2__2__6_ ( .D(n15662), .CK(clk), .Q(template_reg[70])
         );
  QDFFS template_reg_reg_2__2__7_ ( .D(n15661), .CK(clk), .Q(template_reg[71])
         );
  QDFFS cro_mac_reg_0_ ( .D(n13611), .CK(clk), .Q(cro_mac[0]) );
  QDFFS cro_mac_store_reg_0_ ( .D(N7766), .CK(clk), .Q(cro_mac_store[0]) );
  QDFFS cro_mac_reg_1_ ( .D(n13610), .CK(clk), .Q(cro_mac[1]) );
  QDFFS cro_mac_store_reg_1_ ( .D(N7767), .CK(clk), .Q(cro_mac_store[1]) );
  QDFFS cro_mac_reg_2_ ( .D(n13609), .CK(clk), .Q(cro_mac[2]) );
  QDFFS cro_mac_store_reg_2_ ( .D(N7768), .CK(clk), .Q(cro_mac_store[2]) );
  QDFFS cro_mac_reg_3_ ( .D(n13608), .CK(clk), .Q(cro_mac[3]) );
  QDFFS cro_mac_store_reg_3_ ( .D(N7769), .CK(clk), .Q(cro_mac_store[3]) );
  QDFFS cro_mac_reg_4_ ( .D(n13607), .CK(clk), .Q(cro_mac[4]) );
  QDFFS cro_mac_store_reg_4_ ( .D(N7770), .CK(clk), .Q(cro_mac_store[4]) );
  QDFFS cro_mac_reg_5_ ( .D(n13606), .CK(clk), .Q(cro_mac[5]) );
  QDFFS cro_mac_store_reg_5_ ( .D(N7771), .CK(clk), .Q(cro_mac_store[5]) );
  QDFFS cro_mac_reg_6_ ( .D(n13605), .CK(clk), .Q(cro_mac[6]) );
  QDFFS cro_mac_store_reg_6_ ( .D(N7772), .CK(clk), .Q(cro_mac_store[6]) );
  QDFFS cro_mac_reg_7_ ( .D(n13604), .CK(clk), .Q(cro_mac[7]) );
  QDFFS cro_mac_store_reg_7_ ( .D(N7773), .CK(clk), .Q(cro_mac_store[7]) );
  QDFFS cro_mac_reg_8_ ( .D(n13603), .CK(clk), .Q(cro_mac[8]) );
  QDFFS cro_mac_store_reg_8_ ( .D(N7774), .CK(clk), .Q(cro_mac_store[8]) );
  QDFFS cro_mac_reg_9_ ( .D(n13602), .CK(clk), .Q(cro_mac[9]) );
  QDFFS cro_mac_store_reg_9_ ( .D(N7775), .CK(clk), .Q(cro_mac_store[9]) );
  QDFFS cro_mac_reg_10_ ( .D(n13601), .CK(clk), .Q(cro_mac[10]) );
  QDFFS cro_mac_store_reg_10_ ( .D(N7776), .CK(clk), .Q(cro_mac_store[10]) );
  QDFFS cro_mac_reg_11_ ( .D(n13600), .CK(clk), .Q(cro_mac[11]) );
  QDFFS cro_mac_store_reg_11_ ( .D(N7777), .CK(clk), .Q(cro_mac_store[11]) );
  QDFFS cro_mac_reg_12_ ( .D(n13599), .CK(clk), .Q(cro_mac[12]) );
  QDFFS cro_mac_store_reg_12_ ( .D(N7778), .CK(clk), .Q(cro_mac_store[12]) );
  QDFFS cro_mac_reg_13_ ( .D(n13598), .CK(clk), .Q(cro_mac[13]) );
  QDFFS cro_mac_store_reg_13_ ( .D(N7779), .CK(clk), .Q(cro_mac_store[13]) );
  QDFFS cro_mac_reg_14_ ( .D(n13597), .CK(clk), .Q(cro_mac[14]) );
  QDFFS cro_mac_store_reg_14_ ( .D(N7780), .CK(clk), .Q(cro_mac_store[14]) );
  QDFFS cro_mac_reg_15_ ( .D(n13596), .CK(clk), .Q(cro_mac[15]) );
  QDFFS cro_mac_store_reg_15_ ( .D(N7781), .CK(clk), .Q(cro_mac_store[15]) );
  QDFFS cro_mac_reg_16_ ( .D(n13595), .CK(clk), .Q(cro_mac[16]) );
  QDFFS cro_mac_store_reg_16_ ( .D(N7782), .CK(clk), .Q(cro_mac_store[16]) );
  QDFFS cro_mac_reg_17_ ( .D(n13594), .CK(clk), .Q(cro_mac[17]) );
  QDFFS cro_mac_store_reg_17_ ( .D(N7783), .CK(clk), .Q(cro_mac_store[17]) );
  QDFFS cro_mac_reg_18_ ( .D(n13593), .CK(clk), .Q(cro_mac[18]) );
  QDFFS cro_mac_store_reg_18_ ( .D(N7784), .CK(clk), .Q(cro_mac_store[18]) );
  QDFFS cro_mac_reg_19_ ( .D(n13592), .CK(clk), .Q(cro_mac[19]) );
  QDFFS cro_mac_store_reg_19_ ( .D(N7785), .CK(clk), .Q(cro_mac_store[19]) );
  QDFFRBS last_in_valid_reg ( .D(in_valid), .CK(clk), .RB(n15893), .Q(
        last_in_valid) );
  QDFFRBS last_in_valid_d1_reg ( .D(last_in_valid), .CK(clk), .RB(n15893), .Q(
        last_in_valid_d1) );
  QDFFRBS last_in_valid2_reg ( .D(in_valid2), .CK(clk), .RB(n15893), .Q(
        last_in_valid2) );
  QDFFRBS cnt_reg_7_ ( .D(cnt_n[7]), .CK(clk), .RB(n15893), .Q(cnt[7]) );
  QDFFRBS cnt_reg_6_ ( .D(cnt_n[6]), .CK(clk), .RB(n15893), .Q(cnt[6]) );
  QDFFRBS cnt_reg_5_ ( .D(cnt_n[5]), .CK(clk), .RB(n15893), .Q(cnt[5]) );
  QDFFRBS cnt_reg_4_ ( .D(cnt_n[4]), .CK(clk), .RB(n15893), .Q(cnt[4]) );
  QDFFRBS cnt_reg_3_ ( .D(cnt_n[3]), .CK(clk), .RB(n15893), .Q(cnt[3]) );
  QDFFRBS cnt_reg_2_ ( .D(cnt_n[2]), .CK(clk), .RB(n15893), .Q(cnt[2]) );
  QDFFRBS cnt_reg_1_ ( .D(cnt_n[1]), .CK(clk), .RB(n15893), .Q(cnt[1]) );
  QDFFRBS cnt_reg_0_ ( .D(cnt_n[0]), .CK(clk), .RB(n15893), .Q(cnt[0]) );
  QDFFRBS cs_reg_1_ ( .D(n15792), .CK(clk), .RB(n15893), .Q(cs[1]) );
  QDFFRBS cs_d1_reg_1_ ( .D(cs[1]), .CK(clk), .RB(n15893), .Q(cs_d1[1]) );
  QDFFRBS cnt_20_reg_0_ ( .D(cnt_20_n[0]), .CK(clk), .RB(n15893), .Q(cnt_20[0]) );
  QDFFRBS cnt_20_reg_1_ ( .D(cnt_20_n[1]), .CK(clk), .RB(n15893), .Q(cnt_20[1]) );
  QDFFRBS cnt_20_reg_2_ ( .D(cnt_20_n[2]), .CK(clk), .RB(n15893), .Q(cnt_20[2]) );
  QDFFRBS cnt_20_reg_3_ ( .D(cnt_20_n[3]), .CK(clk), .RB(n15893), .Q(cnt_20[3]) );
  QDFFRBS cnt_20_reg_4_ ( .D(cnt_20_n[4]), .CK(clk), .RB(n15893), .Q(cnt_20[4]) );
  QDFFRBS cnt_20_reg_5_ ( .D(cnt_20_n[5]), .CK(clk), .RB(n15893), .Q(cnt_20[5]) );
  QDFFRBS cnt_cro_3_reg_1_ ( .D(n15763), .CK(clk), .RB(n15893), .Q(
        cnt_cro_3[1]) );
  QDFFRBS cnt_cro_y_reg_3_ ( .D(n15745), .CK(clk), .RB(n30454), .Q(
        cnt_cro_y[3]) );
  QDFFRBS cs_reg_2_ ( .D(n15794), .CK(clk), .RB(n30454), .Q(cs[2]) );
  QDFFRBS cs_d1_reg_2_ ( .D(cs[2]), .CK(clk), .RB(n30454), .Q(cs_d1[2]) );
  QDFFRBS cs_reg_0_ ( .D(n15793), .CK(clk), .RB(n30454), .Q(cs[0]) );
  QDFFRBS cs_d1_reg_0_ ( .D(cs[0]), .CK(clk), .RB(n30454), .Q(cs_d1[0]) );
  QDFFRBS action_doing_reg_0_ ( .D(n15760), .CK(clk), .RB(n30454), .Q(
        action_doing[0]) );
  QDFFRBS action_doing_reg_1_ ( .D(n15759), .CK(clk), .RB(n15893), .Q(
        action_doing[1]) );
  QDFFRBS action_doing_reg_2_ ( .D(n15758), .CK(clk), .RB(n15893), .Q(
        action_doing[2]) );
  QDFFRBS cnt_dyn_reg_0_ ( .D(cnt_dyn_n[0]), .CK(clk), .RB(n30454), .Q(
        cnt_dyn[0]) );
  QDFFRBS cnt_dyn_reg_1_ ( .D(n15805), .CK(clk), .RB(n15893), .Q(cnt_dyn[1])
         );
  QDFFRBS cnt_dyn_reg_2_ ( .D(cnt_dyn_n[2]), .CK(clk), .RB(rst_n), .Q(
        cnt_dyn[2]) );
  QDFFRBS cnt_dyn_reg_3_ ( .D(cnt_dyn_n[3]), .CK(clk), .RB(n30454), .Q(
        cnt_dyn[3]) );
  QDFFRBS gray_scale_1_reg_8_ ( .D(gray_scale_1_n[8]), .CK(clk), .RB(n15893), 
        .Q(gray_scale_1[8]) );
  QDFFRBS gray_scale_1_reg_9_ ( .D(gray_scale_1_n[9]), .CK(clk), .RB(rst_n), 
        .Q(gray_scale_1[9]) );
  QDFFRBS gray_scale_2_reg_6_ ( .D(gray_scale_2_n[6]), .CK(clk), .RB(n30454), 
        .Q(gray_scale_2[6]) );
  QDFFRBS gray_scale_2_reg_7_ ( .D(gray_scale_2_n[7]), .CK(clk), .RB(n15893), 
        .Q(gray_scale_2[7]) );
  QDFFRBS gray_scale_0_reg_0_ ( .D(n15744), .CK(clk), .RB(n15893), .Q(
        gray_scale_0[0]) );
  QDFFRBS gray_scale_0_reg_1_ ( .D(n15743), .CK(clk), .RB(n15893), .Q(
        gray_scale_0[1]) );
  QDFFRBS gray_scale_0_reg_2_ ( .D(n15742), .CK(clk), .RB(n15893), .Q(
        gray_scale_0[2]) );
  QDFFRBS gray_scale_0_reg_3_ ( .D(n15741), .CK(clk), .RB(n15893), .Q(
        gray_scale_0[3]) );
  QDFFRBS gray_scale_0_reg_4_ ( .D(n15740), .CK(clk), .RB(n15893), .Q(
        gray_scale_0[4]) );
  QDFFRBS gray_scale_0_reg_5_ ( .D(n15739), .CK(clk), .RB(n15893), .Q(
        gray_scale_0[5]) );
  QDFFRBS gray_scale_0_reg_6_ ( .D(n15738), .CK(clk), .RB(n15893), .Q(
        gray_scale_0[6]) );
  QDFFRBS gray_scale_0_reg_7_ ( .D(n15737), .CK(clk), .RB(n15893), .Q(
        gray_scale_0[7]) );
  QDFFRBS gray_scale_2_reg_0_ ( .D(gray_scale_2_n[0]), .CK(clk), .RB(rst_n), 
        .Q(gray_scale_2[0]) );
  QDFFRBS gray_scale_2_reg_1_ ( .D(gray_scale_2_n[1]), .CK(clk), .RB(rst_n), 
        .Q(gray_scale_2[1]) );
  QDFFRBS gray_scale_2_reg_2_ ( .D(gray_scale_2_n[2]), .CK(clk), .RB(rst_n), 
        .Q(gray_scale_2[2]) );
  QDFFRBS gray_scale_2_reg_3_ ( .D(gray_scale_2_n[3]), .CK(clk), .RB(rst_n), 
        .Q(gray_scale_2[3]) );
  QDFFRBS gray_scale_2_reg_4_ ( .D(gray_scale_2_n[4]), .CK(clk), .RB(n30454), 
        .Q(gray_scale_2[4]) );
  QDFFRBS gray_scale_2_reg_5_ ( .D(gray_scale_2_n[5]), .CK(clk), .RB(n15893), 
        .Q(gray_scale_2[5]) );
  QDFFRBS gray_scale_1_reg_7_ ( .D(n15823), .CK(clk), .RB(n30454), .Q(
        gray_scale_1[7]) );
  QDFFRBS gray_scale_1_reg_6_ ( .D(n15822), .CK(clk), .RB(n15893), .Q(
        gray_scale_1[6]) );
  QDFFRBS gray_scale_1_reg_5_ ( .D(n15821), .CK(clk), .RB(n30454), .Q(
        gray_scale_1[5]) );
  QDFFRBS gray_scale_1_reg_4_ ( .D(n15820), .CK(clk), .RB(n15893), .Q(
        gray_scale_1[4]) );
  QDFFRBS gray_scale_1_reg_3_ ( .D(n15819), .CK(clk), .RB(n30454), .Q(
        gray_scale_1[3]) );
  QDFFRBS gray_scale_1_reg_2_ ( .D(n15818), .CK(clk), .RB(n15893), .Q(
        gray_scale_1[2]) );
  QDFFRBS gray_scale_1_reg_1_ ( .D(n15817), .CK(clk), .RB(n15893), .Q(
        gray_scale_1[1]) );
  QDFFRBS gray_scale_1_reg_0_ ( .D(n15816), .CK(clk), .RB(n15893), .Q(
        gray_scale_1[0]) );
  QDFFRBS cnt_bdyn_reg_8_ ( .D(n15804), .CK(clk), .RB(n15893), .Q(cnt_bdyn[8])
         );
  QDFFRBS cnt_bdyn_reg_7_ ( .D(n15803), .CK(clk), .RB(n15893), .Q(cnt_bdyn[7])
         );
  QDFFRBS cnt_bdyn_reg_6_ ( .D(n15802), .CK(clk), .RB(n15893), .Q(cnt_bdyn[6])
         );
  QDFFRBS cnt_bdyn_reg_5_ ( .D(n15801), .CK(clk), .RB(n15893), .Q(cnt_bdyn[5])
         );
  QDFFRBS cnt_bdyn_reg_4_ ( .D(n15800), .CK(clk), .RB(n15893), .Q(cnt_bdyn[4])
         );
  QDFFRBS mem_we_a_reg_reg ( .D(N442), .CK(clk), .RB(n15893), .Q(mem_we_a_reg)
         );
  QDFFRBS cnt_bdyn_reg_2_ ( .D(n15798), .CK(clk), .RB(n15893), .Q(cnt_bdyn[2])
         );
  QDFFRBS cnt_bdyn_reg_1_ ( .D(n15797), .CK(clk), .RB(n15893), .Q(cnt_bdyn[1])
         );
  QDFFRBS cnt_bdyn_reg_0_ ( .D(n15796), .CK(clk), .RB(n15893), .Q(cnt_bdyn[0])
         );
  QDFFRBS cnt_cro_x_reg_3_ ( .D(n15749), .CK(clk), .RB(n30454), .Q(
        cnt_cro_x[3]) );
  QDFFRBS read_layer_reg_1_ ( .D(n13590), .CK(clk), .RB(n30454), .Q(
        read_layer[1]) );
  QDFFRBS read_layer_reg_0_ ( .D(n13589), .CK(clk), .RB(n15893), .Q(
        read_layer[0]) );
  QDFFRBS set_cnt_reg_0_ ( .D(n13588), .CK(clk), .RB(n15893), .Q(set_cnt[0])
         );
  QDFFRBS set_cnt_reg_1_ ( .D(n13587), .CK(clk), .RB(n15893), .Q(set_cnt[1])
         );
  QDFFRBS set_cnt_reg_2_ ( .D(n13586), .CK(clk), .RB(n15893), .Q(set_cnt[2])
         );
  QDFFRBS out_valid_a1_reg ( .D(n13585), .CK(clk), .RB(n15893), .Q(
        out_valid_a1) );
  QDFFRBS gray_scale_2_s_reg_7_ ( .D(n13584), .CK(clk), .RB(rst_n), .Q(
        gray_scale_2_s[7]) );
  QDFFRBS gray_scale_1_s_reg_0_ ( .D(n13583), .CK(clk), .RB(n15893), .Q(
        gray_scale_1_s[0]) );
  QDFFRBS gray_scale_1_s_reg_1_ ( .D(n13582), .CK(clk), .RB(n15893), .Q(
        gray_scale_1_s[1]) );
  QDFFRBS gray_scale_1_s_reg_2_ ( .D(n13581), .CK(clk), .RB(n30454), .Q(
        gray_scale_1_s[2]) );
  QDFFRBS gray_scale_1_s_reg_3_ ( .D(n13580), .CK(clk), .RB(n30454), .Q(
        gray_scale_1_s[3]) );
  QDFFRBS gray_scale_1_s_reg_4_ ( .D(n13579), .CK(clk), .RB(n30454), .Q(
        gray_scale_1_s[4]) );
  QDFFRBS gray_scale_1_s_reg_5_ ( .D(n13578), .CK(clk), .RB(n15893), .Q(
        gray_scale_1_s[5]) );
  QDFFRBS gray_scale_1_s_reg_6_ ( .D(n13577), .CK(clk), .RB(rst_n), .Q(
        gray_scale_1_s[6]) );
  QDFFRBS gray_scale_1_s_reg_7_ ( .D(n13576), .CK(clk), .RB(n30454), .Q(
        gray_scale_1_s[7]) );
  QDFFRBS gray_scale_0_s_reg_0_ ( .D(n13575), .CK(clk), .RB(n15893), .Q(
        gray_scale_0_s[0]) );
  QDFFRBS gray_scale_0_s_reg_1_ ( .D(n13574), .CK(clk), .RB(n30454), .Q(
        gray_scale_0_s[1]) );
  QDFFRBS gray_scale_0_s_reg_2_ ( .D(n13573), .CK(clk), .RB(n15893), .Q(
        gray_scale_0_s[2]) );
  QDFFRBS gray_scale_0_s_reg_3_ ( .D(n13572), .CK(clk), .RB(n15893), .Q(
        gray_scale_0_s[3]) );
  QDFFRBS gray_scale_0_s_reg_4_ ( .D(n13571), .CK(clk), .RB(n15893), .Q(
        gray_scale_0_s[4]) );
  QDFFRBS gray_scale_0_s_reg_5_ ( .D(n13570), .CK(clk), .RB(n30454), .Q(
        gray_scale_0_s[5]) );
  QDFFRBS gray_scale_0_s_reg_6_ ( .D(n13569), .CK(clk), .RB(n30454), .Q(
        gray_scale_0_s[6]) );
  QDFFRBS gray_scale_0_s_reg_7_ ( .D(n13568), .CK(clk), .RB(n15893), .Q(
        gray_scale_0_s[7]) );
  QDFFRBS gray_scale_2_s_reg_6_ ( .D(n13567), .CK(clk), .RB(n15893), .Q(
        gray_scale_2_s[6]) );
  QDFFRBS gray_scale_2_s_reg_0_ ( .D(n13566), .CK(clk), .RB(n30454), .Q(
        gray_scale_2_s[0]) );
  QDFFRBS gray_scale_2_s_reg_1_ ( .D(n13565), .CK(clk), .RB(n15893), .Q(
        gray_scale_2_s[1]) );
  QDFFRBS gray_scale_2_s_reg_2_ ( .D(n13564), .CK(clk), .RB(n15893), .Q(
        gray_scale_2_s[2]) );
  QDFFRBS gray_scale_2_s_reg_3_ ( .D(n13563), .CK(clk), .RB(n15893), .Q(
        gray_scale_2_s[3]) );
  QDFFRBS gray_scale_2_s_reg_4_ ( .D(n13562), .CK(clk), .RB(n30454), .Q(
        gray_scale_2_s[4]) );
  QDFFRBS gray_scale_2_s_reg_5_ ( .D(n13561), .CK(clk), .RB(n30454), .Q(
        gray_scale_2_s[5]) );
  FA1S DP_OP_989J1_126_3015_U6 ( .A(C1_Z_2), .B(gray_scale_2[2]), .CI(
        DP_OP_989J1_126_3015_n6), .CO(DP_OP_989J1_126_3015_n5), .S(
        C551_DATA2_2) );
  FA1S DP_OP_989J1_126_3015_U4 ( .A(C1_Z_4), .B(gray_scale_2[4]), .CI(
        DP_OP_989J1_126_3015_n4), .CO(DP_OP_989J1_126_3015_n3), .S(
        C551_DATA2_4) );
  FA1S DP_OP_989J1_126_3015_U2 ( .A(C1_Z_6), .B(gray_scale_2[6]), .CI(
        DP_OP_989J1_126_3015_n2), .CO(DP_OP_989J1_126_3015_n1), .S(
        C551_DATA2_6) );
  QDFFRBT cnt_cro_3b3_reg_0_ ( .D(n15761), .CK(clk), .RB(n30454), .Q(
        cnt_cro_3b3[0]) );
  QDFFRBT cnt_cro_3b3_reg_1_ ( .D(n15762), .CK(clk), .RB(n30454), .Q(
        cnt_cro_3b3[1]) );
  QDFFRBS cnt_dyn_base_reg_2_ ( .D(n15754), .CK(clk), .RB(n30454), .Q(
        cnt_dyn_base[2]) );
  QDFFRBN cnt_dyn_base_reg_1_ ( .D(n15789), .CK(clk), .RB(n30454), .Q(
        cnt_dyn_base[1]) );
  QDFFRBP cnt_dyn_base_reg_0_ ( .D(n15755), .CK(clk), .RB(n30454), .Q(
        cnt_dyn_base[0]) );
  QDFFRBS cnt_dyn_base_reg_3_ ( .D(n15753), .CK(clk), .RB(n15893), .Q(
        cnt_dyn_base[3]) );
  QDFFRBS cnt_bdyn_reg_3_ ( .D(n15799), .CK(clk), .RB(n15893), .Q(cnt_bdyn[3])
         );
  QDFFRBS cnt_cro_x_reg_2_ ( .D(n15750), .CK(clk), .RB(n30454), .Q(
        cnt_cro_x[2]) );
  QDFFP medfilt_state_reg_0_ ( .D(n15806), .CK(clk), .Q(medfilt_state[0]) );
  QDFFP medfilt_state_reg_1_ ( .D(N7421), .CK(clk), .Q(medfilt_state[1]) );
  QDFFP medfilt_state_reg_2_ ( .D(N7422), .CK(clk), .Q(medfilt_state[2]) );
  QDFFRBP cnt_cro_x_reg_0_ ( .D(n15752), .CK(clk), .RB(n30454), .Q(
        cnt_cro_x[0]) );
  QDFFRBP cnt_cro_y_reg_0_ ( .D(n15748), .CK(clk), .RB(n15893), .Q(
        cnt_cro_y[0]) );
  QDFFP mem_data_out_reg_shift_1_reg_2__3_ ( .D(mem_data_out_reg_shift_1[11]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[19]) );
  QDFFP medfilt_state_reg_3_ ( .D(n15807), .CK(clk), .Q(medfilt_state[3]) );
  QDFFS medfilt_out_reg_reg_6_ ( .D(n15863), .CK(clk), .Q(medfilt_out_reg[6])
         );
  QDFFS medfilt_out_reg_reg_5_ ( .D(n15862), .CK(clk), .Q(medfilt_out_reg[5])
         );
  QDFFS medfilt_out_reg_reg_4_ ( .D(n15861), .CK(clk), .Q(medfilt_out_reg[4])
         );
  QDFFS medfilt_out_reg_reg_3_ ( .D(n15860), .CK(clk), .Q(medfilt_out_reg[3])
         );
  QDFFS medfilt_out_reg_reg_2_ ( .D(n15859), .CK(clk), .Q(medfilt_out_reg[2])
         );
  FA1 DP_OP_989J1_126_3015_U7 ( .A(C1_Z_1), .B(gray_scale_2[1]), .CI(
        DP_OP_989J1_126_3015_n7), .CO(DP_OP_989J1_126_3015_n6), .S(
        C551_DATA2_1) );
  FA1 DP_OP_989J1_126_3015_U3 ( .A(C1_Z_5), .B(gray_scale_2[5]), .CI(
        DP_OP_989J1_126_3015_n3), .CO(DP_OP_989J1_126_3015_n2), .S(
        C551_DATA2_5) );
  FA1 DP_OP_989J1_126_3015_U5 ( .A(C1_Z_3), .B(gray_scale_2[3]), .CI(
        DP_OP_989J1_126_3015_n5), .CO(DP_OP_989J1_126_3015_n4), .S(
        C551_DATA2_3) );
  QDFFS gray_img_reg_12__0__1_ ( .D(n14340), .CK(clk), .Q(gray_img[1537]) );
  QDFFS gray_img_reg_1__4__1_ ( .D(n14212), .CK(clk), .Q(gray_img[161]) );
  DFFS template_in_reg_reg_3_ ( .D(template[3]), .CK(clk), .Q(
        template_in_reg[3]) );
  DFFS gray_img_reg_6__12__1_ ( .D(n14416), .CK(clk), .Q(gray_img[865]) );
  DFFS gray_img_reg_15__13__0_ ( .D(n13815), .CK(clk), .Q(gray_img[2024]), 
        .QB(intadd_5_B_0_) );
  DFFS gray_img_reg_12__15__0_ ( .D(n13908), .CK(clk), .Q(gray_img[1656]) );
  DFFS gray_img_reg_9__4__1_ ( .D(n14384), .CK(clk), .Q(gray_img[1185]), .QB(
        intadd_83_CI) );
  DFFS gray_img_reg_10__4__1_ ( .D(n14368), .CK(clk), .Q(gray_img[1313]) );
  DFFS gray_img_reg_15__2__1_ ( .D(n14290), .CK(clk), .Q(gray_img[1937]), .QB(
        intadd_151_CI) );
  DFFS gray_img_reg_2__11__0_ ( .D(n14219), .CK(clk), .Q(gray_img[344]) );
  DFFS gray_img_reg_0__14__0_ ( .D(n14260), .CK(clk), .Q(gray_img[112]) );
  DFFS gray_img_reg_7__9__1_ ( .D(n14411), .CK(clk), .Q(gray_img[969]), .QB(
        intadd_98_CI) );
  DFFS gray_img_reg_3__2__1_ ( .D(n14270), .CK(clk), .Q(gray_img[401]), .QB(
        intadd_169_CI) );
  DFFS gray_img_reg_7__1__1_ ( .D(n13686), .CK(clk), .Q(gray_img[905]), .QB(
        intadd_147_CI) );
  DFFS gray_img_reg_2__0__1_ ( .D(n13735), .CK(clk), .Q(gray_img[257]) );
  DFFS mem_data_out_reg_shift_2_reg_1__7_ ( .D(mem_data_out_reg_shift_2[7]), 
        .CK(clk), .Q(mem_data_out_reg_shift_2[15]), .QB(n30455) );
  QDFFRBS out_value_reg ( .D(out_value_a1), .CK(clk), .RB(n30454), .Q(
        out_value) );
  QDFFRBS out_valid_reg ( .D(out_valid_a1), .CK(clk), .RB(n15893), .Q(
        out_valid) );
  QDFFS gray_img_reg_0__5__0_ ( .D(n13809), .CK(clk), .Q(gray_img[40]) );
  QDFFS gray_img_reg_11__8__1_ ( .D(n14348), .CK(clk), .Q(gray_img[1473]) );
  QDFFS gray_img_reg_12__9__1_ ( .D(n14331), .CK(clk), .Q(gray_img[1609]) );
  QDFFS gray_img_reg_2__13__1_ ( .D(n14447), .CK(clk), .Q(gray_img[361]) );
  QDFFS gray_img_reg_7__3__1_ ( .D(n13684), .CK(clk), .Q(gray_img[921]) );
  QDFFS gray_img_reg_9__2__1_ ( .D(n14386), .CK(clk), .Q(gray_img[1169]) );
  QDFFRBN cnt_cro_y_reg_2_ ( .D(n15746), .CK(clk), .RB(n15893), .Q(
        cnt_cro_y[2]) );
  QDFFS gray_img_reg_8__10__1_ ( .D(n14394), .CK(clk), .Q(gray_img[1105]) );
  QDFFS gray_img_reg_10__3__1_ ( .D(n14369), .CK(clk), .Q(gray_img[1305]) );
  QDFFS gray_img_reg_12__13__1_ ( .D(n14327), .CK(clk), .Q(gray_img[1641]) );
  QDFFS gray_img_reg_13__14__1_ ( .D(n14310), .CK(clk), .Q(gray_img[1777]) );
  QDFFS gray_img_reg_10__11__1_ ( .D(n14361), .CK(clk), .Q(gray_img[1369]) );
  QDFFS gray_img_reg_6__15__1_ ( .D(n14413), .CK(clk), .Q(gray_img[889]) );
  QDFFS gray_img_reg_2__10__1_ ( .D(n14450), .CK(clk), .Q(gray_img[337]) );
  QDFFS gray_img_reg_4__4__1_ ( .D(n14036), .CK(clk), .Q(gray_img[545]) );
  QDFFS gray_img_reg_13__1__1_ ( .D(n14323), .CK(clk), .Q(gray_img[1673]) );
  QDFFS gray_img_reg_1__10__1_ ( .D(n14458), .CK(clk), .Q(gray_img[209]) );
  QDFFS gray_img_reg_5__15__1_ ( .D(n14421), .CK(clk), .Q(gray_img[761]) );
  QDFFS gray_img_reg_14__0__1_ ( .D(n14308), .CK(clk), .Q(gray_img[1793]) );
  QDFFS gray_img_reg_9__7__1_ ( .D(n14381), .CK(clk), .Q(gray_img[1209]) );
  QDFFS gray_img_reg_9__6__1_ ( .D(n14382), .CK(clk), .Q(gray_img[1201]) );
  QDFFS gray_img_reg_4__2__1_ ( .D(n14054), .CK(clk), .Q(gray_img[529]) );
  DFFS gray_img_reg_8__15__0_ ( .D(n14075), .CK(clk), .Q(gray_img[1144]) );
  DFFS gray_img_reg_14__15__1_ ( .D(n14293), .CK(clk), .Q(gray_img[1913]) );
  DFFS gray_img_reg_14__15__0_ ( .D(n13844), .CK(clk), .Q(gray_img[1912]) );
  DFFS gray_img_reg_13__15__1_ ( .D(n14309), .CK(clk), .Q(gray_img[1785]), 
        .QB(intadd_32_CI) );
  DFFS gray_img_reg_11__15__1_ ( .D(n14341), .CK(clk), .Q(gray_img[1529]), 
        .QB(intadd_145_CI) );
  DFFS gray_img_reg_1__15__1_ ( .D(n14453), .CK(clk), .Q(gray_img[249]), .QB(
        intadd_123_CI) );
  DFFS gray_img_reg_0__15__1_ ( .D(n14461), .CK(clk), .Q(gray_img[121]) );
  DFFS gray_img_reg_12__12__1_ ( .D(n14328), .CK(clk), .Q(gray_img[1633]), 
        .QB(intadd_36_CI) );
  DFFS gray_img_reg_9__12__1_ ( .D(n14376), .CK(clk), .Q(gray_img[1249]), .QB(
        intadd_72_CI) );
  DFFS gray_img_reg_7__11__1_ ( .D(n14409), .CK(clk), .Q(gray_img[985]) );
  DFFS gray_img_reg_7__10__1_ ( .D(n14410), .CK(clk), .Q(gray_img[977]) );
  DFFS gray_img_reg_6__11__2_ ( .D(n14618), .CK(clk), .Q(gray_img[858]), .QB(
        intadd_96_B_1_) );
  DFFS gray_img_reg_6__11__1_ ( .D(n14417), .CK(clk), .Q(gray_img[857]), .QB(
        intadd_96_CI) );
  DFFS gray_img_reg_6__10__2_ ( .D(n14619), .CK(clk), .Q(gray_img[850]), .QB(
        intadd_97_B_1_) );
  DFFS gray_img_reg_6__10__1_ ( .D(n14418), .CK(clk), .Q(gray_img[849]), .QB(
        intadd_97_CI) );
  DFFS gray_img_reg_4__11__1_ ( .D(n14433), .CK(clk), .Q(gray_img[601]), .QB(
        intadd_106_CI) );
  DFFS gray_img_reg_3__12__1_ ( .D(n14440), .CK(clk), .Q(gray_img[481]), .QB(
        intadd_115_CI) );
  DFFS gray_img_reg_2__12__1_ ( .D(n14448), .CK(clk), .Q(gray_img[353]) );
  DFFS gray_img_reg_1__12__1_ ( .D(n14456), .CK(clk), .Q(gray_img[225]) );
  DFFS gray_img_reg_15__12__1_ ( .D(n14280), .CK(clk), .Q(gray_img[2017]), 
        .QB(intadd_4_CI) );
  DFFS gray_img_reg_3__14__1_ ( .D(n14438), .CK(clk), .Q(gray_img[497]), .QB(
        intadd_112_CI) );
  DFFS gray_img_reg_2__14__1_ ( .D(n14446), .CK(clk), .Q(gray_img[369]) );
  DFFS gray_img_reg_15__14__1_ ( .D(n14278), .CK(clk), .Q(gray_img[2033]), 
        .QB(intadd_1_CI) );
  DFFS gray_img_reg_14__14__0_ ( .D(n13845), .CK(clk), .Q(gray_img[1904]) );
  DFFS gray_img_reg_8__14__1_ ( .D(n14390), .CK(clk), .Q(gray_img[1137]), .QB(
        intadd_69_CI) );
  DFFS gray_img_reg_9__5__1_ ( .D(n14383), .CK(clk), .Q(gray_img[1193]), .QB(
        intadd_82_CI) );
  DFFS gray_img_reg_9__2__2_ ( .D(n14587), .CK(clk), .Q(gray_img[1170]), .QB(
        intadd_85_B_1_) );
  DFFS gray_img_reg_9__0__1_ ( .D(n14388), .CK(clk), .Q(gray_img[1153]), .QB(
        intadd_88_CI) );
  DFFS gray_img_reg_8__5__1_ ( .D(n14399), .CK(clk), .Q(gray_img[1065]) );
  DFFS gray_img_reg_8__5__0_ ( .D(n14085), .CK(clk), .Q(gray_img[1064]) );
  DFFS gray_img_reg_8__1__2_ ( .D(n14604), .CK(clk), .Q(gray_img[1034]), .QB(
        intadd_89_B_1_) );
  DFFS gray_img_reg_8__1__1_ ( .D(n14403), .CK(clk), .Q(gray_img[1033]), .QB(
        intadd_89_CI) );
  DFFS gray_img_reg_3__13__0_ ( .D(n14195), .CK(clk), .Q(gray_img[488]) );
  DFFS gray_img_reg_3__11__1_ ( .D(n14441), .CK(clk), .Q(gray_img[473]), .QB(
        intadd_117_CI) );
  DFFS gray_img_reg_2__11__1_ ( .D(n14449), .CK(clk), .Q(gray_img[345]) );
  DFFS gray_img_reg_0__12__1_ ( .D(n14464), .CK(clk), .Q(gray_img[97]), .QB(
        intadd_125_CI) );
  DFFS gray_img_reg_0__9__1_ ( .D(n14467), .CK(clk), .Q(gray_img[73]), .QB(
        intadd_130_B_0_) );
  DFFS gray_img_reg_7__8__0_ ( .D(n14126), .CK(clk), .Q(gray_img[960]), .QB(
        n30457) );
  DFFS gray_img_reg_3__15__1_ ( .D(n14437), .CK(clk), .Q(gray_img[505]), .QB(
        intadd_111_CI) );
  DFFS gray_img_reg_8__8__0_ ( .D(n14082), .CK(clk), .Q(gray_img[1088]) );
  DFFS gray_img_reg_11__8__0_ ( .D(n13951), .CK(clk), .Q(gray_img[1472]), .QB(
        intadd_186_A_0_) );
  DFFS gray_img_reg_15__8__1_ ( .D(n14284), .CK(clk), .Q(gray_img[1985]), .QB(
        intadd_25_B_0_) );
  DFFS gray_img_reg_15__8__0_ ( .D(n13823), .CK(clk), .Q(gray_img[1984]), .QB(
        intadd_25_A_0_) );
  DFFS gray_img_reg_7__15__1_ ( .D(n14405), .CK(clk), .Q(gray_img[1017]) );
  DFFS gray_img_reg_5__14__1_ ( .D(n14422), .CK(clk), .Q(gray_img[753]), .QB(
        intadd_101_CI) );
  DFFS gray_img_reg_4__14__1_ ( .D(n14430), .CK(clk), .Q(gray_img[625]) );
  DFFS gray_img_reg_9__13__0_ ( .D(n14019), .CK(clk), .Q(gray_img[1256]) );
  DFFS gray_img_reg_15__3__1_ ( .D(n14289), .CK(clk), .Q(gray_img[1945]), .QB(
        intadd_150_CI) );
  DFFS gray_img_reg_14__3__1_ ( .D(n14305), .CK(clk), .Q(gray_img[1817]) );
  DFFS gray_img_reg_8__3__1_ ( .D(n14401), .CK(clk), .Q(gray_img[1049]) );
  DFFS gray_img_reg_9__3__2_ ( .D(n14586), .CK(clk), .Q(gray_img[1178]), .QB(
        intadd_86_B_1_) );
  DFFS gray_img_reg_9__3__1_ ( .D(n14385), .CK(clk), .Q(gray_img[1177]), .QB(
        intadd_86_CI) );
  DFFS gray_img_reg_11__13__1_ ( .D(n14343), .CK(clk), .Q(gray_img[1513]), 
        .QB(intadd_55_CI) );
  DFFS gray_img_reg_9__1__0_ ( .D(n14073), .CK(clk), .Q(gray_img[1160]) );
  DFFS gray_img_reg_10__1__1_ ( .D(n14371), .CK(clk), .Q(gray_img[1289]), .QB(
        intadd_65_CI) );
  DFFS gray_img_reg_9__1__1_ ( .D(n14387), .CK(clk), .Q(gray_img[1161]) );
  DFFS gray_img_reg_9__13__1_ ( .D(n14375), .CK(clk), .Q(gray_img[1257]) );
  DFFS gray_img_reg_8__13__1_ ( .D(n14391), .CK(clk), .Q(gray_img[1129]), .QB(
        intadd_71_CI) );
  DFFS gray_img_reg_9__15__1_ ( .D(n14373), .CK(clk), .Q(gray_img[1273]), .QB(
        intadd_68_CI) );
  DFFS gray_img_reg_9__8__1_ ( .D(n14380), .CK(clk), .Q(gray_img[1217]), .QB(
        intadd_77_CI) );
  DFFS gray_img_reg_8__15__1_ ( .D(n14389), .CK(clk), .Q(gray_img[1145]) );
  DFFS gray_img_reg_8__8__1_ ( .D(n14396), .CK(clk), .Q(gray_img[1089]) );
  DFFS gray_img_reg_13__4__1_ ( .D(n14320), .CK(clk), .Q(gray_img[1697]), .QB(
        intadd_48_CI) );
  DFFS gray_img_reg_15__6__1_ ( .D(n14286), .CK(clk), .Q(gray_img[1969]), .QB(
        intadd_158_CI) );
  DFFS gray_img_reg_14__6__1_ ( .D(n14302), .CK(clk), .Q(gray_img[1841]) );
  DFFS gray_img_reg_13__6__1_ ( .D(n14318), .CK(clk), .Q(gray_img[1713]), .QB(
        intadd_44_CI) );
  DFFS gray_img_reg_11__4__1_ ( .D(n14352), .CK(clk), .Q(gray_img[1441]), .QB(
        intadd_60_CI) );
  DFFS gray_img_reg_11__0__1_ ( .D(n14356), .CK(clk), .Q(gray_img[1409]), .QB(
        intadd_66_CI) );
  DFFS gray_img_reg_10__0__1_ ( .D(n14372), .CK(clk), .Q(gray_img[1281]) );
  DFFS gray_img_reg_15__0__1_ ( .D(n14292), .CK(clk), .Q(gray_img[1921]) );
  DFFS gray_img_reg_13__0__1_ ( .D(n14324), .CK(clk), .Q(gray_img[1665]) );
  DFFS gray_img_reg_13__5__1_ ( .D(n14319), .CK(clk), .Q(gray_img[1705]), .QB(
        intadd_47_CI) );
  DFFS gray_img_reg_11__5__1_ ( .D(n14351), .CK(clk), .Q(gray_img[1449]), .QB(
        intadd_59_CI) );
  DFFS gray_img_reg_10__5__1_ ( .D(n14367), .CK(clk), .Q(gray_img[1321]) );
  DFFS gray_img_reg_11__7__1_ ( .D(n14349), .CK(clk), .Q(gray_img[1465]), .QB(
        intadd_134_CI) );
  DFFS gray_img_reg_13__7__1_ ( .D(n14317), .CK(clk), .Q(gray_img[1721]), .QB(
        intadd_45_CI) );
  DFFS gray_img_reg_10__7__1_ ( .D(n14365), .CK(clk), .Q(gray_img[1337]) );
  DFFS gray_img_reg_14__7__1_ ( .D(n14301), .CK(clk), .Q(gray_img[1849]) );
  DFFS gray_img_reg_15__7__2_ ( .D(n14486), .CK(clk), .Q(gray_img[1978]), .QB(
        intadd_159_B_1_) );
  DFFS gray_img_reg_15__7__1_ ( .D(n14285), .CK(clk), .Q(gray_img[1977]), .QB(
        intadd_159_CI) );
  DFFS gray_img_reg_13__2__1_ ( .D(n14322), .CK(clk), .Q(gray_img[1681]), .QB(
        intadd_50_CI) );
  DFFS gray_img_reg_5__11__1_ ( .D(n14425), .CK(clk), .Q(gray_img[729]) );
  DFFS gray_img_reg_5__9__1_ ( .D(n14427), .CK(clk), .Q(gray_img[713]), .QB(
        intadd_108_CI) );
  DFFS gray_img_reg_0__11__1_ ( .D(n14465), .CK(clk), .Q(gray_img[89]), .QB(
        intadd_188_B_0_) );
  DFFS gray_img_reg_11__10__1_ ( .D(n14346), .CK(clk), .Q(gray_img[1489]) );
  DFFS gray_img_reg_10__10__1_ ( .D(n14362), .CK(clk), .Q(gray_img[1361]), 
        .QB(intadd_140_CI) );
  DFFS gray_img_reg_5__10__1_ ( .D(n14426), .CK(clk), .Q(gray_img[721]) );
  DFFS gray_img_reg_14__12__0_ ( .D(n13847), .CK(clk), .Q(gray_img[1888]) );
  DFFS gray_img_reg_9__12__0_ ( .D(n14020), .CK(clk), .Q(gray_img[1248]), .QB(
        intadd_72_B_0_) );
  DFFS gray_img_reg_7__11__0_ ( .D(n14116), .CK(clk), .Q(gray_img[984]) );
  DFFS gray_img_reg_5__10__0_ ( .D(n14161), .CK(clk), .Q(gray_img[720]) );
  DFFS gray_img_reg_2__10__0_ ( .D(n14220), .CK(clk), .Q(gray_img[336]) );
  DFFS gray_img_reg_13__12__1_ ( .D(n14312), .CK(clk), .Q(gray_img[1761]) );
  DFFS gray_img_reg_3__10__1_ ( .D(n14442), .CK(clk), .Q(gray_img[465]) );
  DFFS gray_img_reg_0__10__1_ ( .D(n14466), .CK(clk), .Q(gray_img[81]) );
  DFFS gray_img_reg_14__8__1_ ( .D(n14300), .CK(clk), .Q(gray_img[1857]) );
  DFFS gray_img_reg_12__8__1_ ( .D(n14332), .CK(clk), .Q(gray_img[1601]), .QB(
        intadd_42_CI) );
  DFFS gray_img_reg_4__15__1_ ( .D(n14429), .CK(clk), .Q(gray_img[633]) );
  DFFS gray_img_reg_4__8__1_ ( .D(n14436), .CK(clk), .Q(gray_img[577]) );
  DFFS gray_img_reg_15__15__1_ ( .D(n14277), .CK(clk), .Q(gray_img[2041]), 
        .QB(intadd_2_A_0_) );
  DFFS gray_img_reg_15__13__1_ ( .D(n14279), .CK(clk), .Q(gray_img[2025]), 
        .QB(intadd_5_CI) );
  DFFS gray_img_reg_10__9__0_ ( .D(n13993), .CK(clk), .Q(gray_img[1352]), .QB(
        n30458) );
  DFFS gray_img_reg_7__10__0_ ( .D(n14117), .CK(clk), .Q(gray_img[976]) );
  DFFS gray_img_reg_0__11__0_ ( .D(n14263), .CK(clk), .Q(gray_img[88]), .QB(
        intadd_188_A_0_) );
  DFFS gray_img_reg_0__10__0_ ( .D(n14264), .CK(clk), .Q(gray_img[80]) );
  DFFS gray_img_reg_0__9__0_ ( .D(n14265), .CK(clk), .Q(gray_img[72]), .QB(
        intadd_130_A_0_) );
  DFFS gray_img_reg_8__7__0_ ( .D(n14083), .CK(clk), .Q(gray_img[1080]) );
  DFFS gray_img_reg_1__14__1_ ( .D(n14454), .CK(clk), .Q(gray_img[241]), .QB(
        intadd_122_CI) );
  DFFS gray_img_reg_0__14__1_ ( .D(n14462), .CK(clk), .Q(gray_img[113]) );
  DFFS gray_img_reg_3__8__2_ ( .D(n14645), .CK(clk), .Q(gray_img[450]), .QB(
        intadd_120_B_1_) );
  DFFS gray_img_reg_3__8__1_ ( .D(n14444), .CK(clk), .Q(gray_img[449]), .QB(
        intadd_120_CI) );
  DFFS gray_img_reg_8__2__1_ ( .D(n14402), .CK(clk), .Q(gray_img[1041]) );
  DFFS gray_img_reg_5__8__1_ ( .D(n14428), .CK(clk), .Q(gray_img[705]), .QB(
        intadd_109_CI) );
  DFFS gray_img_reg_0__8__1_ ( .D(n14468), .CK(clk), .Q(gray_img[65]) );
  DFFS gray_img_reg_0__8__0_ ( .D(n14266), .CK(clk), .Q(gray_img[64]) );
  DFFS gray_img_reg_1__8__1_ ( .D(n14460), .CK(clk), .Q(gray_img[193]), .QB(
        intadd_129_CI) );
  DFFS gray_img_reg_4__13__1_ ( .D(n14431), .CK(clk), .Q(gray_img[617]), .QB(
        intadd_103_CI) );
  DFFS gray_img_reg_6__8__1_ ( .D(n14420), .CK(clk), .Q(gray_img[833]), .QB(
        intadd_99_CI) );
  DFFS gray_img_reg_14__6__0_ ( .D(n13853), .CK(clk), .Q(gray_img[1840]) );
  DFFS gray_img_reg_10__2__0_ ( .D(n14000), .CK(clk), .Q(gray_img[1296]), .QB(
        intadd_62_B_0_) );
  DFFS gray_img_reg_8__3__0_ ( .D(n14087), .CK(clk), .Q(gray_img[1048]) );
  DFFS gray_img_reg_4__10__1_ ( .D(n14434), .CK(clk), .Q(gray_img[593]), .QB(
        intadd_105_CI) );
  DFFS gray_img_reg_1__11__1_ ( .D(n14457), .CK(clk), .Q(gray_img[217]) );
  DFFS gray_img_reg_11__9__1_ ( .D(n14347), .CK(clk), .Q(gray_img[1481]), .QB(
        intadd_57_CI) );
  DFFS gray_img_reg_7__12__1_ ( .D(n14408), .CK(clk), .Q(gray_img[993]), .QB(
        intadd_94_CI) );
  DFFS gray_img_reg_3__9__1_ ( .D(n14443), .CK(clk), .Q(gray_img[457]), .QB(
        intadd_119_CI) );
  DFFS gray_img_reg_15__4__0_ ( .D(n13832), .CK(clk), .Q(gray_img[1952]), .QB(
        intadd_28_A_0_) );
  DFFS gray_img_reg_14__2__1_ ( .D(n14306), .CK(clk), .Q(gray_img[1809]) );
  DFFS gray_img_reg_14__3__0_ ( .D(n13856), .CK(clk), .Q(gray_img[1816]) );
  DFFS gray_img_reg_10__5__0_ ( .D(n13997), .CK(clk), .Q(gray_img[1320]) );
  DFFS gray_img_reg_10__0__0_ ( .D(n14002), .CK(clk), .Q(gray_img[1280]) );
  DFFS gray_img_reg_8__2__0_ ( .D(n14088), .CK(clk), .Q(gray_img[1040]) );
  DFFS gray_img_reg_12__10__0_ ( .D(n13913), .CK(clk), .Q(gray_img[1616]), 
        .QB(intadd_39_B_0_) );
  DFFS gray_img_reg_4__2__2_ ( .D(n14053), .CK(clk), .Q(gray_img[530]), .QB(
        intadd_132_B_1_) );
  DFFS gray_img_reg_4__0__0_ ( .D(n13746), .CK(clk), .Q(gray_img[512]), .QB(
        intadd_8_B_0_) );
  DFFS gray_img_reg_4__0__1_ ( .D(n14072), .CK(clk), .Q(gray_img[513]), .QB(
        intadd_8_CI) );
  DFFS gray_img_reg_6__5__0_ ( .D(n13717), .CK(clk), .Q(gray_img[808]) );
  DFFS gray_img_reg_2__6__0_ ( .D(n13780), .CK(clk), .Q(gray_img[304]), .QB(
        intadd_14_CI) );
  DFFS gray_img_reg_2__6__1_ ( .D(n14150), .CK(clk), .Q(gray_img[305]), .QB(
        intadd_14_B_0_) );
  DFFS gray_img_reg_3__5__1_ ( .D(n14115), .CK(clk), .Q(gray_img[425]) );
  DFFS gray_img_reg_3__3__1_ ( .D(n14269), .CK(clk), .Q(gray_img[409]), .QB(
        intadd_206_CI) );
  DFFS gray_img_reg_5__0__1_ ( .D(n13984), .CK(clk), .Q(gray_img[641]) );
  DFFS gray_img_reg_4__7__0_ ( .D(n13739), .CK(clk), .Q(gray_img[568]), .QB(
        intadd_189_B_0_) );
  DFFS gray_img_reg_4__7__1_ ( .D(n14009), .CK(clk), .Q(gray_img[569]), .QB(
        intadd_189_A_0_) );
  DFFS gray_img_reg_5__4__1_ ( .D(n13699), .CK(clk), .Q(gray_img[673]) );
  DFFS gray_img_reg_7__2__1_ ( .D(n13685), .CK(clk), .Q(gray_img[913]), .QB(
        intadd_156_CI) );
  DFFS gray_img_reg_4__6__1_ ( .D(n14018), .CK(clk), .Q(gray_img[561]) );
  DFFS gray_img_reg_0__0__1_ ( .D(n14276), .CK(clk), .Q(gray_img[1]), .QB(
        intadd_171_B_0_) );
  DFFS gray_img_reg_0__2__1_ ( .D(n13801), .CK(clk), .Q(gray_img[17]), .QB(
        intadd_11_CI) );
  DFFS gray_img_reg_0__2__0_ ( .D(n13802), .CK(clk), .Q(gray_img[16]), .QB(
        intadd_11_B_0_) );
  DFFS gray_img_reg_0__5__1_ ( .D(n14247), .CK(clk), .Q(gray_img[41]), .QB(
        intadd_22_CI) );
  DFFS gray_img_reg_7__0__1_ ( .D(n13687), .CK(clk), .Q(gray_img[897]), .QB(
        intadd_148_CI) );
  DFFS gray_img_reg_1__7__1_ ( .D(n14185), .CK(clk), .Q(gray_img[185]) );
  DFFS gray_img_reg_2__7__1_ ( .D(n14141), .CK(clk), .Q(gray_img[313]), .QB(
        intadd_13_CI) );
  DFFS gray_img_reg_1__7__0_ ( .D(n13793), .CK(clk), .Q(gray_img[184]) );
  DFFS gray_img_reg_2__2__1_ ( .D(n14469), .CK(clk), .Q(gray_img[273]) );
  DFFS gray_img_reg_3__7__1_ ( .D(n14097), .CK(clk), .Q(gray_img[441]) );
  DFFS gray_img_reg_7__5__1_ ( .D(n13682), .CK(clk), .Q(gray_img[937]), .QB(
        intadd_162_CI) );
  DFFS gray_img_reg_4__5__1_ ( .D(n14027), .CK(clk), .Q(gray_img[553]), .QB(
        intadd_137_B_0_) );
  DFFS gray_img_reg_3__7__0_ ( .D(n13763), .CK(clk), .Q(gray_img[440]) );
  DFFS gray_img_reg_3__0__1_ ( .D(n14272), .CK(clk), .Q(gray_img[385]), .QB(
        intadd_153_CI) );
  DFFS gray_img_reg_5__2__1_ ( .D(n13966), .CK(clk), .Q(gray_img[657]) );
  DFFS gray_img_reg_4__5__0_ ( .D(n13741), .CK(clk), .Q(gray_img[552]), .QB(
        intadd_137_A_0_) );
  DFFS gray_img_reg_5__2__0_ ( .D(n13728), .CK(clk), .Q(gray_img[656]) );
  DFFS gray_img_reg_3__1__1_ ( .D(n14271), .CK(clk), .Q(gray_img[393]), .QB(
        intadd_204_CI) );
  DFFS gray_img_reg_5__6__1_ ( .D(n13697), .CK(clk), .Q(gray_img[689]), .QB(
        intadd_142_CI) );
  DFFS gray_img_reg_2__0__0_ ( .D(n13736), .CK(clk), .Q(gray_img[256]) );
  DFFS gray_img_reg_0__6__1_ ( .D(n14238), .CK(clk), .Q(gray_img[49]), .QB(
        intadd_19_B_0_) );
  DFFS gray_img_reg_2__5__1_ ( .D(n14159), .CK(clk), .Q(gray_img[297]), .QB(
        intadd_16_CI) );
  DFFS gray_img_reg_2__5__0_ ( .D(n13781), .CK(clk), .Q(gray_img[296]), .QB(
        intadd_16_B_0_) );
  DFFS medfilt_out_reg_reg_7_ ( .D(n15864), .CK(clk), .Q(medfilt_out_reg[7])
         );
  DFFS template_in_reg_reg_0_ ( .D(template[0]), .CK(clk), .Q(
        template_in_reg[0]) );
  DFFS template_in_reg_reg_1_ ( .D(template[1]), .CK(clk), .Q(
        template_in_reg[1]) );
  DFFS template_in_reg_reg_2_ ( .D(template[2]), .CK(clk), .Q(
        template_in_reg[2]) );
  DFFS template_in_reg_reg_4_ ( .D(template[4]), .CK(clk), .Q(
        template_in_reg[4]) );
  DFFS template_in_reg_reg_5_ ( .D(template[5]), .CK(clk), .Q(
        template_in_reg[5]) );
  DFFS template_in_reg_reg_6_ ( .D(template[6]), .CK(clk), .Q(
        template_in_reg[6]) );
  DFFS template_in_reg_reg_7_ ( .D(template[7]), .CK(clk), .Q(
        template_in_reg[7]) );
  HA1S DP_OP_989J1_126_3015_U8 ( .A(C1_Z_0), .B(gray_scale_2[0]), .C(
        DP_OP_989J1_126_3015_n7), .S(C551_DATA2_0) );
  DFFS mem_data_out_reg_shift_1_reg_2__5_ ( .D(mem_data_out_reg_shift_1[13]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[21]), .QB(n30456) );
  QDFFN mem_data_out_reg_shift_1_reg_2__4_ ( .D(mem_data_out_reg_shift_1[12]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[20]) );
  QDFFN mem_data_out_reg_shift_1_reg_2__2_ ( .D(mem_data_out_reg_shift_1[10]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[18]) );
  QDFFN mem_data_out_reg_shift_1_reg_2__1_ ( .D(mem_data_out_reg_shift_1[9]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[17]) );
  QDFFN mem_data_out_reg_shift_1_reg_2__7_ ( .D(mem_data_out_reg_shift_1[15]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[23]) );
  QDFFN mem_data_out_reg_shift_1_reg_2__6_ ( .D(mem_data_out_reg_shift_1[14]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[22]) );
  QDFFN mem_data_out_reg_shift_1_reg_2__0_ ( .D(mem_data_out_reg_shift_1[8]), 
        .CK(clk), .Q(mem_data_out_reg_shift_1[16]) );
  QDFFRBP cnt_cro_y_reg_1_ ( .D(n15747), .CK(clk), .RB(n30454), .Q(
        cnt_cro_y[1]) );
  QDFFRBN cnt_cro_x_reg_1_ ( .D(n15751), .CK(clk), .RB(n30454), .Q(
        cnt_cro_x[1]) );
  QDFFRBN cnt_cro_3_reg_0_ ( .D(n15764), .CK(clk), .RB(n30454), .Q(
        cnt_cro_3[0]) );
  NR2 U15941 ( .I1(n29680), .I2(n26207), .O(n26327) );
  NR2 U15942 ( .I1(n29680), .I2(n26650), .O(n29739) );
  NR2 U15943 ( .I1(n29680), .I2(n27928), .O(n28136) );
  NR2 U15944 ( .I1(n29680), .I2(n28643), .O(n28706) );
  NR2 U15945 ( .I1(n29680), .I2(n25548), .O(n25604) );
  INV1S U15946 ( .I(n19092), .O(n29734) );
  FA1S U15947 ( .A(n30417), .B(gray_scale_0[3]), .CI(n23050), .CO(n23051) );
  INV1S U15948 ( .I(n19127), .O(n18734) );
  NR2 U15949 ( .I1(n24772), .I2(n24771), .O(n24870) );
  ND3 U15950 ( .I1(n24522), .I2(n24521), .I3(n24520), .O(n24819) );
  BUF1 U15951 ( .I(n22945), .O(n15915) );
  BUF1 U15952 ( .I(n22769), .O(n15918) );
  FA1S U15953 ( .A(n17169), .B(n17168), .CI(n17167), .CO(n17962), .S(n17366)
         );
  ND2P U15954 ( .I1(n24759), .I2(n24420), .O(n24758) );
  NR2T U15955 ( .I1(n15987), .I2(n24255), .O(n24514) );
  INV2 U15956 ( .I(n18450), .O(n25315) );
  ND3 U15957 ( .I1(n23942), .I2(n23941), .I3(n23940), .O(n24480) );
  BUF2 U15958 ( .I(n16119), .O(n15914) );
  BUF2 U15959 ( .I(n16150), .O(n15913) );
  BUF2 U15960 ( .I(n16156), .O(n15909) );
  BUF2 U15961 ( .I(n16296), .O(n15902) );
  BUF2 U15962 ( .I(n16500), .O(n15900) );
  INV3 U15963 ( .I(n15867), .O(n15895) );
  INV3 U15964 ( .I(n15947), .O(n15876) );
  MOAI1S U15965 ( .A1(n24380), .A2(n24660), .B1(n24379), .B2(n24658), .O(
        n24352) );
  INV3 U15966 ( .I(n16363), .O(n15872) );
  INV3 U15967 ( .I(n15910), .O(n15911) );
  BUF2 U15968 ( .I(n24639), .O(n24698) );
  OR2 U15969 ( .I1(n16211), .I2(n16203), .O(n16518) );
  ND2P U15970 ( .I1(n16140), .I2(n16138), .O(n17505) );
  ND2P U15971 ( .I1(n16141), .I2(n16140), .O(n17381) );
  ND2P U15972 ( .I1(n16140), .I2(n16122), .O(n17704) );
  OR2 U15973 ( .I1(n16125), .I2(n16159), .O(n16210) );
  INV1S U15974 ( .I(n16142), .O(n15907) );
  INV1S U15975 ( .I(n16134), .O(n15910) );
  OR2P U15976 ( .I1(n16147), .I2(n16136), .O(n16209) );
  OR2P U15977 ( .I1(n16136), .I2(n16135), .O(n16203) );
  INV3 U15978 ( .I(n16147), .O(n16135) );
  OAI12HS U15979 ( .B1(n23712), .B2(n23711), .A1(n23710), .O(n23735) );
  XOR2HS U15980 ( .I1(n16102), .I2(n16101), .O(n16154) );
  XNR2HS U15981 ( .I1(n16110), .I2(n16109), .O(n16148) );
  INV3 U15982 ( .I(n23949), .O(n23896) );
  OAI12HS U15983 ( .B1(n23906), .B2(n24292), .A1(n23717), .O(n24294) );
  NR2P U15984 ( .I1(n23666), .I2(n23650), .O(n24316) );
  INV1S U15985 ( .I(n24273), .O(n24613) );
  ND3 U15986 ( .I1(n23774), .I2(n23773), .I3(n23772), .O(n24607) );
  OAI12HS U15987 ( .B1(n23781), .B2(n24327), .A1(n23780), .O(n24579) );
  ND3 U15988 ( .I1(n23787), .I2(n23786), .I3(n23785), .O(n24578) );
  ND3 U15989 ( .I1(n23754), .I2(n23753), .I3(n23752), .O(n24557) );
  AN2 U15990 ( .I1(n24919), .I2(n30242), .O(n23781) );
  NR2P U15991 ( .I1(n23991), .I2(n23990), .O(n24646) );
  NR2P U15992 ( .I1(n24013), .I2(n24012), .O(n24638) );
  AN4B1S U15993 ( .I1(n17284), .I2(n17283), .I3(n17282), .B1(n17281), .O(
        n17307) );
  ND3S U15994 ( .I1(n16222), .I2(n16221), .I3(n16220), .O(n16291) );
  ND3S U15995 ( .I1(n16737), .I2(n16736), .I3(n16735), .O(n16783) );
  BUF2 U15996 ( .I(n17521), .O(n15912) );
  INV3 U15997 ( .I(n15946), .O(n15898) );
  INV1S U15998 ( .I(n24754), .O(n24665) );
  OAI12HS U15999 ( .B1(n24137), .B2(n24136), .A1(n24135), .O(n24203) );
  FA1S U16000 ( .A(cro_mac[11]), .B(n17959), .CI(n17958), .CO(n17979), .S(
        n17961) );
  NR2P U16001 ( .I1(n24263), .I2(n24614), .O(n23961) );
  NR2P U16002 ( .I1(cnt_cro_3b3[1]), .I2(n16111), .O(n16113) );
  ND3S U16003 ( .I1(n24202), .I2(n24201), .I3(n24200), .O(n24477) );
  MOAI1S U16004 ( .A1(n30413), .A2(n30409), .B1(n16006), .B2(action_done), .O(
        n16007) );
  OA112 U16005 ( .C1(n24620), .C2(n24619), .A1(n24618), .B1(n24617), .O(n24801) );
  AN2 U16006 ( .I1(action_doing[2]), .I2(n30410), .O(n16006) );
  NR2 U16007 ( .I1(n30384), .I2(n16007), .O(n16047) );
  NR3H U16008 ( .I1(medfilt_state[0]), .I2(medfilt_state[2]), .I3(n23637), .O(
        n18464) );
  ND3S U16009 ( .I1(cs[2]), .I2(n16089), .I3(n18145), .O(n30384) );
  ND2P U16010 ( .I1(n16011), .I2(n16047), .O(n25374) );
  INV1S U16011 ( .I(n24755), .O(n24868) );
  NR2 U16012 ( .I1(n29680), .I2(n23240), .O(n28806) );
  NR2 U16013 ( .I1(n29680), .I2(n28180), .O(n28247) );
  NR2 U16014 ( .I1(n29680), .I2(n28517), .O(n28671) );
  NR2 U16015 ( .I1(n29680), .I2(n26797), .O(n27355) );
  HA1 U16016 ( .A(image[0]), .B(gray_scale_1[0]), .C(n30347), .S(n30350) );
  INV3 U16017 ( .I(n29734), .O(n15888) );
  INV3CK U16018 ( .I(n29837), .O(n28530) );
  NR2 U16019 ( .I1(n29680), .I2(n18092), .O(n29350) );
  BUF1CK U16020 ( .I(n22809), .O(n15921) );
  BUF1CK U16021 ( .I(n22827), .O(n15919) );
  NR2P U16022 ( .I1(n16210), .I2(n16204), .O(n15866) );
  OR2 U16023 ( .I1(n16205), .I2(n16196), .O(n15867) );
  ND2 U16024 ( .I1(n16047), .I2(n16006), .O(n16048) );
  INV4 U16025 ( .I(n16048), .O(n27447) );
  INV3 U16026 ( .I(n16048), .O(n15889) );
  OR2 U16027 ( .I1(n16208), .I2(n16209), .O(n15868) );
  INV3 U16028 ( .I(n15940), .O(n15901) );
  AN2 U16029 ( .I1(n25315), .I2(n27222), .O(n15869) );
  BUF1S U16030 ( .I(n27314), .O(n15925) );
  BUF1CK U16031 ( .I(n15924), .O(n15887) );
  BUF1S U16032 ( .I(n15924), .O(n15926) );
  BUF1CK U16033 ( .I(n15924), .O(n15881) );
  BUF1CK U16034 ( .I(n27314), .O(n15880) );
  INV1S U16035 ( .I(n29843), .O(n27314) );
  BUF1S U16036 ( .I(n27314), .O(n15924) );
  INV1S U16037 ( .I(n29849), .O(n30057) );
  BUF1CK U16038 ( .I(n15936), .O(n15883) );
  BUF1S U16039 ( .I(n30057), .O(n15934) );
  BUF1S U16040 ( .I(n15934), .O(n15938) );
  BUF1CK U16041 ( .I(n15934), .O(n15882) );
  BUF1S U16042 ( .I(n15934), .O(n15935) );
  BUF1S U16043 ( .I(n30057), .O(n15936) );
  BUF1S U16044 ( .I(n15934), .O(n15939) );
  BUF1CK U16045 ( .I(n15936), .O(n15937) );
  BUF1S U16046 ( .I(n15930), .O(n15933) );
  BUF1S U16047 ( .I(n27512), .O(n15928) );
  BUF1CK U16048 ( .I(n15930), .O(n15884) );
  BUF1S U16049 ( .I(n15928), .O(n15929) );
  BUF1S U16050 ( .I(n15930), .O(n15932) );
  BUF1CK U16051 ( .I(n15929), .O(n15886) );
  INV1S U16052 ( .I(n29884), .O(n27512) );
  BUF1S U16053 ( .I(n27512), .O(n15930) );
  BUF1CK U16054 ( .I(n15930), .O(n15885) );
  BUF1S U16055 ( .I(n15930), .O(n15931) );
  AN2 U16056 ( .I1(n17556), .I2(n17555), .O(n15870) );
  AN2 U16057 ( .I1(n16590), .I2(n16589), .O(n15871) );
  NR2 U16058 ( .I1(n29680), .I2(n26569), .O(n29579) );
  NR2 U16059 ( .I1(n29680), .I2(n29822), .O(n29880) );
  NR2 U16060 ( .I1(n29680), .I2(n26692), .O(n30020) );
  OR2 U16061 ( .I1(n29680), .I2(n23534), .O(n28585) );
  NR2 U16062 ( .I1(n29680), .I2(n23623), .O(n26931) );
  OR2 U16063 ( .I1(n29680), .I2(n25815), .O(n25933) );
  OR2 U16064 ( .I1(n29680), .I2(n16044), .O(n26846) );
  OR2 U16065 ( .I1(n29680), .I2(n28395), .O(n28597) );
  OR2 U16066 ( .I1(n29680), .I2(n29940), .O(n30001) );
  OR2 U16067 ( .I1(n29680), .I2(n26411), .O(n26470) );
  OR2 U16068 ( .I1(n29680), .I2(n26611), .O(n29477) );
  NR2 U16069 ( .I1(n29680), .I2(n29232), .O(n29273) );
  OR2 U16070 ( .I1(n29680), .I2(n28889), .O(n28947) );
  OR2 U16071 ( .I1(n29680), .I2(n29639), .O(n30099) );
  OR2 U16072 ( .I1(n29680), .I2(n27593), .O(n27698) );
  INV3 U16073 ( .I(n15869), .O(n29680) );
  INV4 U16074 ( .I(n17505), .O(n17744) );
  BUF4 U16075 ( .I(n16301), .O(n15873) );
  INV3 U16076 ( .I(n16379), .O(n15874) );
  INV2 U16077 ( .I(n15868), .O(n15875) );
  ND2 U16078 ( .I1(n20988), .I2(n25374), .O(n28452) );
  ND2 U16079 ( .I1(n20982), .I2(n25374), .O(n28601) );
  ND2 U16080 ( .I1(n21047), .I2(n25374), .O(n28208) );
  ND2 U16081 ( .I1(n20994), .I2(n25374), .O(n28943) );
  ND2 U16082 ( .I1(n18140), .I2(n25374), .O(n30121) );
  ND2 U16083 ( .I1(n21000), .I2(n25374), .O(n29186) );
  ND2 U16084 ( .I1(n21035), .I2(n25374), .O(n28121) );
  ND2 U16085 ( .I1(n25327), .I2(n25374), .O(n30032) );
  INV3 U16086 ( .I(n16518), .O(n15877) );
  ND2 U16087 ( .I1(n25375), .I2(n25374), .O(n27834) );
  INV4 U16088 ( .I(n15944), .O(n15878) );
  ND2 U16089 ( .I1(n23412), .I2(n25374), .O(n26932) );
  BUF3 U16090 ( .I(n16325), .O(n15879) );
  ND2 U16091 ( .I1(n21041), .I2(n25374), .O(n27702) );
  ND2 U16092 ( .I1(n21018), .I2(n25374), .O(n30006) );
  ND2 U16093 ( .I1(n21053), .I2(n25374), .O(n27814) );
  ND2 U16094 ( .I1(n21023), .I2(n25374), .O(n27685) );
  ND2 U16095 ( .I1(n21071), .I2(n25374), .O(n30070) );
  ND2 U16096 ( .I1(n21029), .I2(n25374), .O(n27779) );
  ND2 U16097 ( .I1(n20912), .I2(n25374), .O(n29598) );
  ND2 U16098 ( .I1(n16055), .I2(n25374), .O(n26842) );
  OR2 U16099 ( .I1(n30424), .I2(n30419), .O(n30420) );
  BUF1 U16100 ( .I(n27314), .O(n15927) );
  NR2P U16101 ( .I1(n16120), .I2(n16159), .O(n16126) );
  ND2 U16102 ( .I1(medfilt_cnt_d1[0]), .I2(n18641), .O(n24996) );
  INV2 U16103 ( .I(n29825), .O(n15890) );
  INV2 U16104 ( .I(n29831), .O(n15891) );
  INV2 U16105 ( .I(n25291), .O(n15892) );
  ND2 U16106 ( .I1(mem_data_a_out[0]), .I2(n16010), .O(n18733) );
  NR2P U16107 ( .I1(n21157), .I2(n21144), .O(n22664) );
  NR2P U16108 ( .I1(n21144), .I2(n21147), .O(n22863) );
  AN2 U16109 ( .I1(n19127), .I2(medfilt_out_reg[7]), .O(n19128) );
  ND2 U16110 ( .I1(n18139), .I2(n18138), .O(n24999) );
  ND2 U16111 ( .I1(n18470), .I2(n16053), .O(n18543) );
  ND2 U16112 ( .I1(n18095), .I2(n16054), .O(n18510) );
  ND2 U16113 ( .I1(medfilt_cnt2_d1[0]), .I2(n16050), .O(n18537) );
  ND2 U16114 ( .I1(medfilt_cnt2_d1[1]), .I2(n16051), .O(n18571) );
  ND2 U16115 ( .I1(n18094), .I2(n16051), .O(n18509) );
  ND2 U16116 ( .I1(n18469), .I2(n16050), .O(n18542) );
  ND2 U16117 ( .I1(medfilt_cnt_d1[2]), .I2(n18137), .O(n25050) );
  ND2 U16118 ( .I1(cnt_bdyn_d1[0]), .I2(n16053), .O(n18538) );
  ND2 U16119 ( .I1(cnt_bdyn_d1[1]), .I2(n16054), .O(n18572) );
  ND2 U16120 ( .I1(n18137), .I2(n18136), .O(n24997) );
  ND2 U16121 ( .I1(cnt_dyn_d1[1]), .I2(n18138), .O(n24973) );
  BUF2 U16122 ( .I(rst_n), .O(n15893) );
  ND2S U16123 ( .I1(n18002), .I2(n18001), .O(n18012) );
  ND2S U16124 ( .I1(n18048), .I2(n18047), .O(n18052) );
  OA12 U16125 ( .B1(n30199), .B2(n30203), .A1(n30200), .O(n30197) );
  ND3 U16126 ( .I1(n24191), .I2(n24190), .I3(n24189), .O(n24500) );
  INV2 U16127 ( .I(n16786), .O(n17873) );
  BUF4CK U16128 ( .I(n24199), .O(n15922) );
  OR2 U16129 ( .I1(n29680), .I2(n25689), .O(n25740) );
  OR2 U16130 ( .I1(n29680), .I2(n28325), .O(n28456) );
  AN4B1S U16131 ( .I1(n16563), .I2(n16562), .I3(n16561), .B1(n16560), .O(
        n16586) );
  INV4 U16132 ( .I(n15907), .O(n15908) );
  OR2 U16133 ( .I1(n27447), .I2(n20323), .O(n20586) );
  OR2 U16134 ( .I1(n27447), .I2(n20335), .O(n20354) );
  INV4 U16135 ( .I(n15866), .O(n15894) );
  BUF3 U16136 ( .I(n16129), .O(n17765) );
  OR2 U16137 ( .I1(n27447), .I2(n18626), .O(n20296) );
  OR2 U16138 ( .I1(n27447), .I2(n18487), .O(n20477) );
  OR2 U16139 ( .I1(n27447), .I2(n18674), .O(n20833) );
  OR2 U16140 ( .I1(n27447), .I2(n18611), .O(n20159) );
  OR2 U16141 ( .I1(n27447), .I2(n18861), .O(n20392) );
  OR2 U16142 ( .I1(n27447), .I2(n18775), .O(n20836) );
  OR2 U16143 ( .I1(n27447), .I2(n18705), .O(n20427) );
  OR2 U16144 ( .I1(n27447), .I2(n18479), .O(n20541) );
  OR2 U16145 ( .I1(n27447), .I2(n18830), .O(n20517) );
  OR2 U16146 ( .I1(n27447), .I2(n18484), .O(n20522) );
  ND2 U16147 ( .I1(n19667), .I2(n30005), .O(n20435) );
  OR2 U16148 ( .I1(n27447), .I2(n18760), .O(n20395) );
  OR2 U16149 ( .I1(n27447), .I2(n18568), .O(n20843) );
  ND2 U16150 ( .I1(n19807), .I2(n30005), .O(n20480) );
  OR2 U16151 ( .I1(n27447), .I2(n18888), .O(n20362) );
  OR2 U16152 ( .I1(n27447), .I2(n18954), .O(n20449) );
  OR2 U16153 ( .I1(n27447), .I2(n18816), .O(n20512) );
  OR2 U16154 ( .I1(n27447), .I2(n18742), .O(n20430) );
  OR2 U16155 ( .I1(n27447), .I2(n18690), .O(n20849) );
  OR2 U16156 ( .I1(n27447), .I2(n18651), .O(n20486) );
  OR2 U16157 ( .I1(n27447), .I2(n18683), .O(n20846) );
  OR2 U16158 ( .I1(n27447), .I2(n18504), .O(n20379) );
  OR2 U16159 ( .I1(n27447), .I2(n18521), .O(n20824) );
  OR2 U16160 ( .I1(n27447), .I2(n18596), .O(n20129) );
  OR2 U16161 ( .I1(n27447), .I2(n18896), .O(n20602) );
  OR2 U16162 ( .I1(n27447), .I2(n18790), .O(n20547) );
  OR2 U16163 ( .I1(n27447), .I2(n18708), .O(n20550) );
  OR2 U16164 ( .I1(n27447), .I2(n18923), .O(n20591) );
  OR2 U16165 ( .I1(n27447), .I2(n18663), .O(n20839) );
  OR2 U16166 ( .I1(n27447), .I2(n18848), .O(n20376) );
  OR2 U16167 ( .I1(n27447), .I2(n18965), .O(n20719) );
  OR2 U16168 ( .I1(n27447), .I2(n18936), .O(n20209) );
  OR2 U16169 ( .I1(n27447), .I2(n18608), .O(n19970) );
  OR2 U16170 ( .I1(n27447), .I2(n18693), .O(n20472) );
  OR2 U16171 ( .I1(n27447), .I2(n18988), .O(n20734) );
  OR2 U16172 ( .I1(n27447), .I2(n18586), .O(n20725) );
  OR2 U16173 ( .I1(n27447), .I2(n18752), .O(n20202) );
  OR2 U16174 ( .I1(n27447), .I2(n20866), .O(n20881) );
  ND2 U16175 ( .I1(n19846), .I2(n30005), .O(n20617) );
  OR2 U16176 ( .I1(n27447), .I2(n18813), .O(n20319) );
  OR2 U16177 ( .I1(n27447), .I2(n18836), .O(n20731) );
  OR2 U16178 ( .I1(n27447), .I2(n18985), .O(n19955) );
  OR2 U16179 ( .I1(n27447), .I2(n18855), .O(n20746) );
  OR2 U16180 ( .I1(n27447), .I2(n19002), .O(n20702) );
  OR2 U16181 ( .I1(n27447), .I2(n18899), .O(n20389) );
  OR2 U16182 ( .I1(n27447), .I2(n18768), .O(n20655) );
  OR2 U16183 ( .I1(n27447), .I2(n18980), .O(n20528) );
  OR2 U16184 ( .I1(n27447), .I2(n18605), .O(n20596) );
  OR2 U16185 ( .I1(n27447), .I2(n18823), .O(n20695) );
  ND2 U16186 ( .I1(n19731), .I2(n30005), .O(n20757) );
  OR2 U16187 ( .I1(n27447), .I2(n18809), .O(n20424) );
  OR2 U16188 ( .I1(n27447), .I2(n18968), .O(n20722) );
  OR2 U16189 ( .I1(n27447), .I2(n18878), .O(n20373) );
  OR2 U16190 ( .I1(n27447), .I2(n18736), .O(n20556) );
  OR2 U16191 ( .I1(n27447), .I2(n18833), .O(n20737) );
  OR2 U16192 ( .I1(n27447), .I2(n18669), .O(n20857) );
  ND2 U16193 ( .I1(n19415), .I2(n30005), .O(n20235) );
  OR2 U16194 ( .I1(n27447), .I2(n18602), .O(n20599) );
  ND2 U16195 ( .I1(n25943), .I2(n30005), .O(n25942) );
  ND2 U16196 ( .I1(n19408), .I2(n30005), .O(n20614) );
  OR2 U16197 ( .I1(n27447), .I2(n18589), .O(n20124) );
  OR2 U16198 ( .I1(n27447), .I2(n18739), .O(n20142) );
  OR2 U16199 ( .I1(n27447), .I2(n18702), .O(n20035) );
  OR2 U16200 ( .I1(n27447), .I2(n18677), .O(n20854) );
  OR2 U16201 ( .I1(n27447), .I2(n18549), .O(n20054) );
  OR2 U16202 ( .I1(n27447), .I2(n18957), .O(n20728) );
  OR2 U16203 ( .I1(n27447), .I2(n18599), .O(n20293) );
  ND2 U16204 ( .I1(n19688), .I2(n30005), .O(n20311) );
  ND2 U16205 ( .I1(n19891), .I2(n30005), .O(n20631) );
  OR2 U16206 ( .I1(n27447), .I2(n18960), .O(n20463) );
  ND2 U16207 ( .I1(n19726), .I2(n30005), .O(n20760) );
  OR2 U16208 ( .I1(n27447), .I2(n18910), .O(n20384) );
  OR2 U16209 ( .I1(n27447), .I2(n18826), .O(n20709) );
  OR2 U16210 ( .I1(n27447), .I2(n18666), .O(n20821) );
  OR2 U16211 ( .I1(n27447), .I2(n18885), .O(n20193) );
  OR2 U16212 ( .I1(n27447), .I2(n18995), .O(n20743) );
  OR2 U16213 ( .I1(n27447), .I2(n18926), .O(n20147) );
  OR2 U16214 ( .I1(n27447), .I2(n18893), .O(n20605) );
  OR2 U16215 ( .I1(n27447), .I2(n18713), .O(n20531) );
  OR2 U16216 ( .I1(n27447), .I2(n18492), .O(n20525) );
  OR2 U16217 ( .I1(n27447), .I2(n18977), .O(n20504) );
  OR2 U16218 ( .I1(n27447), .I2(n18539), .O(n20562) );
  OR2 U16219 ( .I1(n27447), .I2(n18648), .O(n20568) );
  OR2 U16220 ( .I1(n27447), .I2(n18680), .O(n20862) );
  OR2 U16221 ( .I1(n27447), .I2(n18660), .O(n20099) );
  ND2 U16222 ( .I1(n19789), .I2(n30005), .O(n20608) );
  OR2 U16223 ( .I1(n27447), .I2(n18544), .O(n20559) );
  OR2 U16224 ( .I1(n27447), .I2(n18747), .O(n20571) );
  OR2 U16225 ( .I1(n27447), .I2(n18904), .O(n20212) );
  OR2 U16226 ( .I1(n27447), .I2(n18757), .O(n20827) );
  OR2 U16227 ( .I1(n27447), .I2(n18495), .O(n20063) );
  OR2 U16228 ( .I1(n27447), .I2(n18616), .O(n20184) );
  OR2 U16229 ( .I1(n27447), .I2(n18654), .O(n20452) );
  NR2 U16230 ( .I1(n16198), .I2(n16196), .O(n16119) );
  ND2 U16231 ( .I1(n19833), .I2(n30005), .O(n20274) );
  OR2 U16232 ( .I1(n27447), .I2(n18851), .O(n20740) );
  ND2 U16233 ( .I1(n19759), .I2(n30005), .O(n20316) );
  OR2 U16234 ( .I1(n27447), .I2(n18686), .O(n20496) );
  OR2 U16235 ( .I1(n27447), .I2(n18471), .O(n20156) );
  OR2 U16236 ( .I1(n27447), .I2(n18511), .O(n20368) );
  OR2 U16237 ( .I1(n27447), .I2(n18718), .O(n20553) );
  OR2 U16238 ( .I1(n27447), .I2(n18643), .O(n20082) );
  OR2 U16239 ( .I1(n27447), .I2(n18573), .O(n20811) );
  OR2 U16240 ( .I1(n27447), .I2(n18534), .O(n20534) );
  OR2 U16241 ( .I1(n27447), .I2(n18516), .O(n20787) );
  OR2 U16242 ( .I1(n27447), .I2(n18998), .O(n20684) );
  OR2 U16243 ( .I1(n27447), .I2(n18951), .O(n20544) );
  INV2 U16244 ( .I(n15868), .O(n15896) );
  ND2 U16245 ( .I1(n19800), .I2(n30005), .O(n20491) );
  OR2 U16246 ( .I1(n27447), .I2(n18845), .O(n20583) );
  ND2 U16247 ( .I1(n19773), .I2(n30005), .O(n20255) );
  OR2 U16248 ( .I1(n27447), .I2(n18763), .O(n20509) );
  ND2 U16249 ( .I1(n19699), .I2(n30005), .O(n20240) );
  OR2 U16250 ( .I1(n27447), .I2(n18771), .O(n20814) );
  OR2 U16251 ( .I1(n27447), .I2(n18929), .O(n20580) );
  OR2 U16252 ( .I1(n27447), .I2(n18974), .O(n20440) );
  ND2 U16253 ( .I1(n19826), .I2(n30005), .O(n20620) );
  OR2 U16254 ( .I1(n27447), .I2(n18778), .O(n20716) );
  OR2 U16255 ( .I1(n27447), .I2(n18907), .O(n20365) );
  OR2 U16256 ( .I1(n27447), .I2(n18657), .O(n20565) );
  ND2 U16257 ( .I1(n19664), .I2(n30005), .O(n20611) );
  OR2 U16258 ( .I1(n27447), .I2(n18858), .O(n20359) );
  BUF3 U16259 ( .I(n17716), .O(n15897) );
  BUF2 U16260 ( .I(n16368), .O(n15899) );
  OR2S U16261 ( .I1(n16060), .I2(n16046), .O(n16041) );
  OR2S U16262 ( .I1(n27667), .I2(n27669), .O(n27584) );
  INV3 U16263 ( .I(n16495), .O(n15903) );
  INV2 U16264 ( .I(n27447), .O(n15904) );
  ND3 U16265 ( .I1(cnt_dyn_d1[0]), .I2(cnt_dyn_d1[3]), .I3(n18642), .O(n24998)
         );
  OR2 U16266 ( .I1(n24997), .I2(n24996), .O(n25366) );
  ND3 U16267 ( .I1(cnt_dyn_d1[3]), .I2(n18642), .I3(n18478), .O(n25051) );
  OR2 U16268 ( .I1(n25050), .I2(n25049), .O(n25341) );
  MAO222S U16269 ( .A1(n26200), .B1(gray_img[742]), .C1(n26172), .O(n26173) );
  INV3 U16270 ( .I(n15889), .O(n30005) );
  OR2 U16271 ( .I1(n24972), .I2(n25049), .O(n25357) );
  OR2 U16272 ( .I1(n24972), .I2(n24996), .O(n25352) );
  ND2 U16273 ( .I1(cnt_dyn_d1[0]), .I2(n16052), .O(n18821) );
  BUF1 U16274 ( .I(n15889), .O(n28534) );
  ND2 U16275 ( .I1(n16049), .I2(n18477), .O(n18883) );
  ND2 U16276 ( .I1(medfilt_cnt_d1[0]), .I2(n16049), .O(n18819) );
  ND2 U16277 ( .I1(n18641), .I2(n18477), .O(n25049) );
  ND3P U16278 ( .I1(n23770), .I2(n23769), .I3(n23768), .O(n24599) );
  AOI12H U16279 ( .B1(mem_data_a_out[6]), .B2(n16010), .A1(n18097), .O(n29825)
         );
  AOI12H U16280 ( .B1(mem_data_a_out[5]), .B2(n16010), .A1(n18518), .O(n29831)
         );
  NR2P U16281 ( .I1(n30452), .I2(n30361), .O(n22679) );
  AOI12HP U16282 ( .B1(mem_data_a_out[7]), .B2(n16010), .A1(n19128), .O(n25291) );
  NR2P U16283 ( .I1(n30251), .I2(n30308), .O(n21137) );
  ND3 U16284 ( .I1(n30367), .I2(n30393), .I3(n30130), .O(n30131) );
  INV1 U16285 ( .I(n22889), .O(n22797) );
  NR2P U16286 ( .I1(n21151), .I2(n21156), .O(n21089) );
  INV2 U16287 ( .I(n22383), .O(n15905) );
  NR2P U16288 ( .I1(n21157), .I2(n21131), .O(n22686) );
  NR2P U16289 ( .I1(n30411), .I2(n30380), .O(n30226) );
  NR2P U16290 ( .I1(n21154), .I2(n21156), .O(n21090) );
  NR2P U16291 ( .I1(n21159), .I2(n30306), .O(n21155) );
  NR2P U16292 ( .I1(n21151), .I2(n21153), .O(n21152) );
  NR2P U16293 ( .I1(n21145), .I2(n21146), .O(n22934) );
  NR2P U16294 ( .I1(n21154), .I2(n21157), .O(n21096) );
  NR2P U16295 ( .I1(n21154), .I2(n21146), .O(n21120) );
  NR2P U16296 ( .I1(n21131), .I2(n21147), .O(n22513) );
  NR2P U16297 ( .I1(n18167), .I2(n18181), .O(n18165) );
  NR2P U16298 ( .I1(n18181), .I2(n18180), .O(n18182) );
  NR2P U16299 ( .I1(n21131), .I2(n21156), .O(n22610) );
  NR2P U16300 ( .I1(n21154), .I2(n30306), .O(n22935) );
  NR2P U16301 ( .I1(n18178), .I2(n18177), .O(n18179) );
  NR2P U16302 ( .I1(action_doing[2]), .I2(n25315), .O(n16010) );
  NR2P U16303 ( .I1(n18173), .I2(n18156), .O(n18157) );
  NR2P U16304 ( .I1(n21131), .I2(n21146), .O(n22625) );
  NR2P U16305 ( .I1(n18178), .I2(n18181), .O(n18161) );
  NR2P U16306 ( .I1(n21157), .I2(n21145), .O(n21106) );
  NR2P U16307 ( .I1(n18167), .I2(n18177), .O(n18155) );
  NR2P U16308 ( .I1(n21159), .I2(n21156), .O(n22936) );
  NR2P U16309 ( .I1(n21158), .I2(n21145), .O(n22770) );
  OR2 U16310 ( .I1(n18571), .I2(n18566), .O(n25287) );
  NR2P U16311 ( .I1(n18175), .I2(n18167), .O(n18168) );
  OR2 U16312 ( .I1(n18532), .I2(n18566), .O(n25054) );
  OR2 U16313 ( .I1(n18577), .I2(n18566), .O(n25066) );
  NR2P U16314 ( .I1(n18173), .I2(n18180), .O(n18169) );
  NR2P U16315 ( .I1(n21153), .I2(n21131), .O(n22630) );
  NR2P U16316 ( .I1(n18167), .I2(n18173), .O(n18158) );
  NR2P U16317 ( .I1(n18175), .I2(n18178), .O(n18159) );
  INV3 U16318 ( .I(n18464), .O(n24118) );
  NR2P U16319 ( .I1(n18178), .I2(n18173), .O(n18174) );
  NR2P U16320 ( .I1(n21153), .I2(n21145), .O(n21097) );
  OR2 U16321 ( .I1(n18532), .I2(n18576), .O(n25058) );
  NR2P U16322 ( .I1(n21145), .I2(n30306), .O(n22703) );
  OR2 U16323 ( .I1(n18571), .I2(n18576), .O(n25293) );
  OR2 U16324 ( .I1(cnt_cro_3[1]), .I2(n16103), .O(n16226) );
  ND3 U16325 ( .I1(n30413), .I2(action_doing[1]), .I3(action_doing[0]), .O(
        n18450) );
  ND2 U16326 ( .I1(cnt_dyn_d1[2]), .I2(n18139), .O(n25052) );
  NR2P U16327 ( .I1(n30388), .I2(n18400), .O(n18401) );
  NR2P U16328 ( .I1(n17576), .I2(n17577), .O(n18007) );
  ND3 U16329 ( .I1(n24492), .I2(n24491), .I3(n24490), .O(n24817) );
  NR2F U16330 ( .I1(n24325), .I2(n24263), .O(n24262) );
  ND2 U16331 ( .I1(n30451), .I2(n30330), .O(n21138) );
  ND3 U16332 ( .I1(n24386), .I2(n24385), .I3(n24384), .O(n24387) );
  AOI12H U16333 ( .B1(n17923), .B2(n30170), .A1(n17922), .O(n17972) );
  BUF2 U16334 ( .I(n23662), .O(n15906) );
  NR2P U16335 ( .I1(n24476), .I2(n24475), .O(n24888) );
  NR2 U16336 ( .I1(n16164), .I2(n16196), .O(n16142) );
  ND3 U16337 ( .I1(n24643), .I2(n24642), .I3(n24641), .O(n24749) );
  AOI22S U16338 ( .A1(n16000), .A2(gray_img[1124]), .B1(n17751), .B2(
        gray_img[1636]), .O(n16909) );
  INV3 U16339 ( .I(n16003), .O(n17786) );
  NR2 U16340 ( .I1(n16212), .I2(n16174), .O(n16156) );
  NR2 U16341 ( .I1(n16168), .I2(n16196), .O(n16134) );
  INV3 U16342 ( .I(n24849), .O(n24850) );
  NR2P U16343 ( .I1(n24424), .I2(n24423), .O(n24853) );
  INV1S U16344 ( .I(n16461), .O(n17521) );
  OR2 U16345 ( .I1(n16208), .I2(n16207), .O(n16477) );
  ND3 U16346 ( .I1(n24261), .I2(n24260), .I3(n24259), .O(n24851) );
  OAI112H U16347 ( .C1(n24785), .C2(n24868), .A1(n24784), .B1(n24783), .O(
        n24883) );
  INV3 U16348 ( .I(n16002), .O(n17779) );
  NR2 U16349 ( .I1(n16205), .I2(n16173), .O(n16150) );
  OAI112H U16350 ( .C1(n24801), .C2(n24868), .A1(n24800), .B1(n24799), .O(
        n24816) );
  OR2 U16351 ( .I1(n23807), .I2(n23905), .O(n23717) );
  INV2 U16352 ( .I(n16127), .O(n15916) );
  INV4 U16353 ( .I(n15916), .O(n15917) );
  NR2 U16354 ( .I1(n16213), .I2(n16168), .O(n16127) );
  OR2 U16355 ( .I1(n16208), .I2(n16196), .O(n16363) );
  ND3 U16356 ( .I1(n24467), .I2(n24873), .I3(n24825), .O(n24469) );
  ND3 U16357 ( .I1(n24451), .I2(n24450), .I3(n24449), .O(n24825) );
  NR2T U16358 ( .I1(n23738), .I2(n23735), .O(n24325) );
  OR2P U16359 ( .I1(n16152), .I2(n16151), .O(n16174) );
  INV2 U16360 ( .I(n22896), .O(n22540) );
  BUF2 U16361 ( .I(n23665), .O(n15920) );
  INV1 U16362 ( .I(n17197), .O(n16265) );
  NR2P U16363 ( .I1(n24674), .I2(n24676), .O(n24060) );
  NR2T U16364 ( .I1(n24039), .I2(n24038), .O(n24674) );
  NR2 U16365 ( .I1(n23951), .I2(n24600), .O(n23884) );
  INV2 U16366 ( .I(n24598), .O(n23951) );
  NR2T U16367 ( .I1(n16168), .I2(n16203), .O(n16137) );
  ND2P U16368 ( .I1(n16126), .I2(n16158), .O(n16168) );
  AOI12H U16369 ( .B1(n23798), .B2(n23797), .A1(n23796), .O(n23799) );
  INV2 U16370 ( .I(n24320), .O(n24582) );
  BUF2 U16371 ( .I(n24453), .O(n15923) );
  NR2P U16372 ( .I1(n24341), .I2(n23680), .O(n23681) );
  NR2 U16373 ( .I1(n24600), .I2(n23950), .O(n23795) );
  NR2 U16374 ( .I1(n24542), .I2(n24280), .O(n23763) );
  OAI12H U16375 ( .B1(n23781), .B2(n24283), .A1(n23742), .O(n24542) );
  OAI12H U16376 ( .B1(mem_data_out_reg_shift_1[22]), .B2(n23677), .A1(n23676), 
        .O(n23680) );
  INV2 U16377 ( .I(mem_data_out_reg_shift_1[20]), .O(n24327) );
  ND2S U16378 ( .I1(n24918), .I2(mem_data_out_reg_shift_0[20]), .O(n23780) );
  ND3P U16379 ( .I1(n23749), .I2(n23748), .I3(n23747), .O(n24546) );
  FA1 U16380 ( .A(image[5]), .B(gray_scale_1[5]), .CI(n30339), .CO(n30336), 
        .S(n30340) );
  FA1 U16381 ( .A(image[4]), .B(gray_scale_1[4]), .CI(n30341), .CO(n30339), 
        .S(n30342) );
  OAI12H U16382 ( .B1(n23890), .B2(n23889), .A1(n23888), .O(n23949) );
  NR2P U16383 ( .I1(n24589), .I2(n24315), .O(n23792) );
  ND2 U16384 ( .I1(n24315), .I2(n24589), .O(n23790) );
  ND2S U16385 ( .I1(n24589), .I2(n24592), .O(n23879) );
  NR2 U16386 ( .I1(n24592), .I2(n24589), .O(n23881) );
  ND2 U16387 ( .I1(n23966), .I2(n24589), .O(n23969) );
  OAI12H U16388 ( .B1(n23781), .B2(n30456), .A1(n23776), .O(n24589) );
  INV2 U16389 ( .I(n24312), .O(n24592) );
  NR2P U16390 ( .I1(n23895), .I2(n24427), .O(n24764) );
  INV2 U16391 ( .I(n23891), .O(n23895) );
  NR2P U16392 ( .I1(n24444), .I2(n24443), .O(n24873) );
  INV2 U16393 ( .I(n24607), .O(n24276) );
  ND3P U16394 ( .I1(n23758), .I2(n23757), .I3(n23756), .O(n24856) );
  MOAI1H U16395 ( .A1(n24052), .A2(n24051), .B1(mem_data_out_reg_shift_1[22]), 
        .B2(n24050), .O(n24345) );
  MOAI1 U16396 ( .A1(n15983), .A2(n23675), .B1(n24268), .B2(
        mem_data_out_reg_shift_1[22]), .O(n23676) );
  INV2 U16397 ( .I(n24599), .O(n23950) );
  ND2T U16398 ( .I1(n24842), .I2(n24843), .O(n24896) );
  FA1 U16399 ( .A(image[7]), .B(gray_scale_1[7]), .CI(n30285), .CO(n30287), 
        .S(n18055) );
  FA1 U16400 ( .A(image[6]), .B(gray_scale_1[6]), .CI(n30336), .CO(n30285), 
        .S(n30337) );
  MAOI1 U16401 ( .A1(n30288), .A2(gray_scale_1[9]), .B1(n30288), .B2(
        gray_scale_1[9]), .O(n30289) );
  HA1P U16402 ( .A(gray_scale_1[8]), .B(n30287), .C(n30288), .S(n30286) );
  AN3S U16403 ( .I1(n23659), .I2(n23658), .I3(n23657), .O(n15983) );
  AOI12HS U16404 ( .B1(n24098), .B2(n24097), .A1(n24096), .O(n24137) );
  NR2 U16405 ( .I1(n24158), .I2(n24157), .O(n24159) );
  MAO222S U16406 ( .A1(n24138), .B1(n24196), .C1(n24141), .O(n24158) );
  NR2P U16407 ( .I1(n24156), .I2(n24155), .O(n24157) );
  OAI12H U16408 ( .B1(n24066), .B2(n24065), .A1(n24064), .O(n24169) );
  AOI12HS U16409 ( .B1(n24021), .B2(n24020), .A1(n24019), .O(n24066) );
  OR2S U16410 ( .I1(n24245), .I2(n24486), .O(n24249) );
  MAO222 U16411 ( .A1(n22969), .B1(gray_img[967]), .C1(n22968), .O(n22994) );
  MAO222 U16412 ( .A1(n22971), .B1(gray_img[966]), .C1(n22967), .O(n22968) );
  MAO222 U16413 ( .A1(n22966), .B1(gray_img[965]), .C1(n22965), .O(n22967) );
  MAO222S U16414 ( .A1(n22982), .B1(gray_img[847]), .C1(n22981), .O(n23295) );
  MAO222 U16415 ( .A1(n22980), .B1(gray_img[846]), .C1(n22979), .O(n22981) );
  MAO222 U16416 ( .A1(n27175), .B1(gray_img[845]), .C1(n22978), .O(n22979) );
  MAO222 U16417 ( .A1(n22977), .B1(gray_img[844]), .C1(n22976), .O(n22978) );
  MAO222 U16418 ( .A1(n25027), .B1(n25028), .C1(n23238), .O(n23239) );
  MAO222 U16419 ( .A1(n25762), .B1(n25766), .C1(n23237), .O(n23238) );
  MAO222 U16420 ( .A1(n28685), .B1(n28689), .C1(n23236), .O(n23237) );
  MAO222 U16421 ( .A1(n28690), .B1(n28694), .C1(n23235), .O(n23236) );
  MAO222S U16422 ( .A1(n25319), .B1(n25320), .C1(n18132), .O(n18133) );
  MAO222 U16423 ( .A1(n18135), .B1(n18144), .C1(n18131), .O(n18132) );
  MAO222 U16424 ( .A1(n30043), .B1(n30041), .C1(n18130), .O(n18131) );
  MAO222 U16425 ( .A1(n30049), .B1(n30047), .C1(n18129), .O(n18130) );
  MAO222S U16426 ( .A1(n27885), .B1(n27884), .C1(n27883), .O(n27886) );
  MAO222 U16427 ( .A1(n27888), .B1(n27892), .C1(n27882), .O(n27883) );
  MAO222 U16428 ( .A1(n28824), .B1(n28822), .C1(n27881), .O(n27882) );
  MAO222 U16429 ( .A1(n28829), .B1(n28827), .C1(n27880), .O(n27881) );
  MAO222S U16430 ( .A1(n27734), .B1(gray_img[183]), .C1(n27733), .O(n27786) );
  MAO222 U16431 ( .A1(n27730), .B1(gray_img[181]), .C1(n27729), .O(n27731) );
  MAO222 U16432 ( .A1(n27721), .B1(gray_img[191]), .C1(n27720), .O(n27735) );
  MAO222 U16433 ( .A1(n27719), .B1(gray_img[190]), .C1(n27718), .O(n27720) );
  MAO222 U16434 ( .A1(n27717), .B1(gray_img[189]), .C1(n27716), .O(n27718) );
  MAO222 U16435 ( .A1(n27715), .B1(gray_img[188]), .C1(n27714), .O(n27716) );
  MAO222S U16436 ( .A1(n25007), .B1(n25008), .C1(n23579), .O(n23580) );
  MAO222 U16437 ( .A1(n25637), .B1(n25635), .C1(n23578), .O(n23579) );
  MAO222 U16438 ( .A1(n25724), .B1(n25722), .C1(n23577), .O(n23578) );
  MAO222 U16439 ( .A1(n25729), .B1(n25727), .C1(n23576), .O(n23577) );
  MAO222S U16440 ( .A1(n23159), .B1(n23158), .C1(n23157), .O(n23160) );
  MAO222 U16441 ( .A1(n23188), .B1(n23192), .C1(n23156), .O(n23157) );
  MAO222 U16442 ( .A1(n23183), .B1(n23187), .C1(n23155), .O(n23156) );
  MAO222S U16443 ( .A1(n23178), .B1(n23182), .C1(n23154), .O(n23155) );
  MAO222 U16444 ( .A1(n27926), .B1(n27925), .C1(n27924), .O(n27927) );
  MAO222 U16445 ( .A1(n27929), .B1(n27933), .C1(n27923), .O(n27924) );
  MAO222 U16446 ( .A1(n27934), .B1(n27938), .C1(n27922), .O(n27923) );
  MAO222S U16447 ( .A1(n27939), .B1(n27943), .C1(n27921), .O(n27922) );
  MAO222S U16448 ( .A1(n25206), .B1(n25207), .C1(n23533), .O(n23534) );
  MOAI1S U16449 ( .A1(n23532), .A2(n23531), .B1(n23544), .B2(n23548), .O(
        n23533) );
  MAO222 U16450 ( .A1(n23332), .B1(n23331), .C1(n23330), .O(n23333) );
  MAO222 U16451 ( .A1(n23350), .B1(n23354), .C1(n23329), .O(n23330) );
  MAO222 U16452 ( .A1(n23340), .B1(n23344), .C1(n23328), .O(n23329) );
  MAO222 U16453 ( .A1(n23355), .B1(n23359), .C1(n23327), .O(n23328) );
  MAO222 U16454 ( .A1(n26367), .B1(n26366), .C1(n26365), .O(n26368) );
  MAO222 U16455 ( .A1(n26370), .B1(n26374), .C1(n26364), .O(n26365) );
  MAO222 U16456 ( .A1(n26450), .B1(n26448), .C1(n26363), .O(n26364) );
  MOAI1S U16457 ( .A1(n26362), .A2(n26361), .B1(n26453), .B2(n26455), .O(
        n26363) );
  MAO222 U16458 ( .A1(n26174), .B1(gray_img[743]), .C1(n26173), .O(n26198) );
  MAO222S U16459 ( .A1(n26171), .B1(gray_img[741]), .C1(n26170), .O(n26172) );
  MAO222 U16460 ( .A1(n27037), .B1(gray_img[735]), .C1(n27036), .O(n27106) );
  MAO222 U16461 ( .A1(n27035), .B1(gray_img[734]), .C1(n27034), .O(n27036) );
  MAO222 U16462 ( .A1(n27025), .B1(gray_img[727]), .C1(n27024), .O(n27038) );
  MAO222S U16463 ( .A1(n27023), .B1(gray_img[726]), .C1(n27022), .O(n27024) );
  MAO222S U16464 ( .A1(n27021), .B1(gray_img[725]), .C1(n27020), .O(n27022) );
  MAO222S U16465 ( .A1(n27019), .B1(gray_img[724]), .C1(n27018), .O(n27020) );
  MAO222S U16466 ( .A1(n25249), .B1(n25250), .C1(n23407), .O(n23408) );
  MAO222S U16467 ( .A1(n26867), .B1(n26865), .C1(n23406), .O(n23407) );
  MAO222 U16468 ( .A1(n26908), .B1(n26906), .C1(n23405), .O(n23406) );
  MAO222 U16469 ( .A1(n26913), .B1(n26911), .C1(n23404), .O(n23405) );
  MAO222S U16470 ( .A1(n27580), .B1(gray_img[119]), .C1(n27579), .O(n27586) );
  MAO222S U16471 ( .A1(n27578), .B1(gray_img[118]), .C1(n27577), .O(n27579) );
  MAO222S U16472 ( .A1(n27576), .B1(gray_img[117]), .C1(n27575), .O(n27577) );
  MAO222 U16473 ( .A1(n27568), .B1(gray_img[127]), .C1(n27567), .O(n27699) );
  MAO222 U16474 ( .A1(n27566), .B1(gray_img[126]), .C1(n27565), .O(n27567) );
  MAO222 U16475 ( .A1(n27564), .B1(gray_img[125]), .C1(n27563), .O(n27565) );
  MAO222S U16476 ( .A1(n27562), .B1(gray_img[124]), .C1(n27561), .O(n27563) );
  ND2S U16477 ( .I1(action_doing[1]), .I2(action_doing[2]), .O(n18458) );
  MUX2S U16478 ( .A(gray_img[1289]), .B(gray_img[1417]), .S(n29991), .O(n29706) );
  MUX2S U16479 ( .A(gray_img[953]), .B(gray_img[825]), .S(n28725), .O(n28241)
         );
  MUX2S U16480 ( .A(n29597), .B(n26322), .S(gray_img[304]), .O(n26323) );
  MUX2S U16481 ( .A(n15904), .B(n29740), .S(gray_img[512]), .O(n29733) );
  MUX2S U16482 ( .A(gray_img[1217]), .B(gray_img[1089]), .S(n28669), .O(n28589) );
  MUX2S U16483 ( .A(n30044), .B(n26842), .S(gray_img[40]), .O(n23485) );
  MUX2S U16484 ( .A(n30056), .B(n28840), .S(gray_img[136]), .O(n28816) );
  MUX2S U16485 ( .A(n15904), .B(n28728), .S(gray_img[408]), .O(n28729) );
  MUX2S U16486 ( .A(n29566), .B(n25751), .S(gray_img[928]), .O(n23585) );
  MUX2S U16487 ( .A(n30056), .B(n30121), .S(gray_img[128]), .O(n23362) );
  MUX2S U16488 ( .A(n29587), .B(n30021), .S(gray_img[912]), .O(n30022) );
  MUX2S U16489 ( .A(n30044), .B(n29481), .S(gray_img[768]), .O(n29483) );
  MUX2S U16490 ( .A(n15904), .B(n28248), .S(gray_img[280]), .O(n28217) );
  MUX2S U16491 ( .A(n30005), .B(n28137), .S(gray_img[696]), .O(n28138) );
  MUX2S U16492 ( .A(n15904), .B(n28707), .S(gray_img[272]), .O(n28681) );
  MUX2S U16493 ( .A(n15904), .B(n29994), .S(gray_img[640]), .O(n29995) );
  MUX2S U16494 ( .A(n15904), .B(n28672), .S(gray_img[544]), .O(n28673) );
  MUX2S U16495 ( .A(n29597), .B(n27845), .S(gray_img[152]), .O(n27847) );
  MUX2S U16496 ( .A(n30005), .B(n27702), .S(gray_img[56]), .O(n27704) );
  MUX2S U16497 ( .A(n30050), .B(n26924), .S(gray_img[32]), .O(n23627) );
  MUX2S U16498 ( .A(n30044), .B(n26842), .S(gray_img[43]), .O(n16067) );
  MUX2S U16499 ( .A(n29566), .B(n29344), .S(gray_img[668]), .O(n23204) );
  ND2S U16500 ( .I1(n28530), .I2(n29344), .O(n23203) );
  AN4B1S U16501 ( .I1(n17083), .I2(n17082), .I3(n17081), .B1(n17080), .O(
        n17090) );
  ND2S U16502 ( .I1(n25037), .I2(cnt_cro_3b3[1]), .O(n16100) );
  ND2S U16503 ( .I1(n24578), .I2(n24582), .O(n23850) );
  AO12S U16504 ( .B1(n23914), .B2(mem_data_out_reg_shift_1[17]), .A1(
        mem_data_out_reg_shift_1[16]), .O(n23647) );
  NR2 U16505 ( .I1(n24131), .I2(n24123), .O(n24134) );
  AN4B1S U16506 ( .I1(n17045), .I2(n17044), .I3(n17043), .B1(n17042), .O(
        n17068) );
  ND2S U16507 ( .I1(n16591), .I2(cnt_cro_3b3[0]), .O(n16594) );
  AO222S U16508 ( .A1(template_reg[36]), .A2(n17581), .B1(template_reg[44]), 
        .B2(n17580), .C1(n17579), .C2(template_reg[28]), .O(n16591) );
  AN2S U16509 ( .I1(n24859), .I2(n24856), .O(n15981) );
  NR2P U16510 ( .I1(n23795), .I2(n23775), .O(n23798) );
  MAO222S U16511 ( .A1(gray_img[1233]), .B1(gray_img[1232]), .C1(n28302), .O(
        n28303) );
  NR2 U16512 ( .I1(n24283), .I2(n23672), .O(n23654) );
  NR2 U16513 ( .I1(n24327), .I2(n23672), .O(n23656) );
  OR2S U16514 ( .I1(n23826), .I2(n23905), .O(n23723) );
  ND2S U16515 ( .I1(n16597), .I2(cnt_cro_3b3[0]), .O(n16600) );
  AO222S U16516 ( .A1(template_reg[39]), .A2(n17581), .B1(template_reg[47]), 
        .B2(n17580), .C1(n17579), .C2(template_reg[31]), .O(n16597) );
  AO222S U16517 ( .A1(template_reg[14]), .A2(n17581), .B1(template_reg[6]), 
        .B2(n17579), .C1(n17580), .C2(template_reg[22]), .O(n16792) );
  ND3S U16518 ( .I1(n16790), .I2(n16789), .I3(n16788), .O(n16791) );
  AO222S U16519 ( .A1(template_reg[13]), .A2(n17581), .B1(template_reg[5]), 
        .B2(n17579), .C1(n17580), .C2(template_reg[21]), .O(n16980) );
  AO222S U16520 ( .A1(template_reg[35]), .A2(n17581), .B1(template_reg[43]), 
        .B2(n17580), .C1(n17579), .C2(template_reg[27]), .O(n16397) );
  AO222S U16521 ( .A1(template_reg[33]), .A2(n17581), .B1(template_reg[41]), 
        .B2(n17580), .C1(n17579), .C2(template_reg[25]), .O(n17358) );
  NR2P U16522 ( .I1(n23956), .I2(n23681), .O(n23682) );
  MAO222S U16523 ( .A1(n23222), .B1(gray_img[802]), .C1(n23221), .O(n23223) );
  MAO222S U16524 ( .A1(gray_img[800]), .B1(gray_img[801]), .C1(n23220), .O(
        n23221) );
  MAO222S U16525 ( .A1(n29618), .B1(gray_img[770]), .C1(n29617), .O(n29619) );
  MAO222S U16526 ( .A1(gray_img[768]), .B1(gray_img[769]), .C1(intadd_148_CI), 
        .O(n29617) );
  MAO222S U16527 ( .A1(n26956), .B1(gray_img[169]), .C1(intadd_22_CI), .O(
        n26957) );
  MAO222S U16528 ( .A1(n29276), .B1(gray_img[794]), .C1(n29275), .O(n29277) );
  MAO222S U16529 ( .A1(gray_img[793]), .B1(gray_img[792]), .C1(n29274), .O(
        n29275) );
  MAO222S U16530 ( .A1(n23140), .B1(gray_img[1842]), .C1(n23139), .O(n23141)
         );
  MAO222S U16531 ( .A1(gray_img[1840]), .B1(gray_img[1841]), .C1(intadd_158_CI), .O(n23139) );
  MAO222S U16532 ( .A1(n25998), .B1(gray_img[1650]), .C1(n25997), .O(n25999)
         );
  MAO222S U16533 ( .A1(gray_img[1648]), .B1(gray_img[1649]), .C1(n25996), .O(
        n25997) );
  MAO222S U16534 ( .A1(n27894), .B1(gray_img[1402]), .C1(n27893), .O(n27895)
         );
  MAO222S U16535 ( .A1(gray_img[1401]), .B1(gray_img[1400]), .C1(intadd_145_CI), .O(n27893) );
  MAO222S U16536 ( .A1(gray_img[1346]), .B1(n23502), .C1(n23501), .O(n23503)
         );
  MAO222S U16537 ( .A1(n23500), .B1(intadd_186_A_0_), .C1(gray_img[1345]), .O(
        n23501) );
  MAO222S U16538 ( .A1(n23301), .B1(gray_img[1266]), .C1(n23300), .O(n23302)
         );
  MAO222S U16539 ( .A1(gray_img[1265]), .B1(gray_img[1264]), .C1(intadd_69_CI), 
        .O(n23300) );
  MAO222S U16540 ( .A1(n28855), .B1(gray_img[1082]), .C1(n28854), .O(n28856)
         );
  MAO222S U16541 ( .A1(gray_img[1081]), .B1(gray_img[1080]), .C1(n28853), .O(
        n28854) );
  MAO222S U16542 ( .A1(n23022), .B1(gray_img[1066]), .C1(n23021), .O(n23023)
         );
  MAO222S U16543 ( .A1(gray_img[1065]), .B1(gray_img[1064]), .C1(intadd_82_CI), 
        .O(n23021) );
  MAO222S U16544 ( .A1(gray_img[1041]), .B1(gray_img[1040]), .C1(n29800), .O(
        n29801) );
  MAO222S U16545 ( .A1(n26390), .B1(gray_img[1018]), .C1(n26389), .O(n26391)
         );
  MAO222S U16546 ( .A1(gray_img[1017]), .B1(gray_img[1016]), .C1(n26388), .O(
        n26389) );
  MAO222S U16547 ( .A1(n26334), .B1(gray_img[634]), .C1(n26333), .O(n26335) );
  MAO222S U16548 ( .A1(gray_img[633]), .B1(gray_img[632]), .C1(n26332), .O(
        n26333) );
  MAO222S U16549 ( .A1(n27612), .B1(gray_img[378]), .C1(n27611), .O(n27613) );
  MAO222S U16550 ( .A1(gray_img[376]), .B1(gray_img[377]), .C1(intadd_111_CI), 
        .O(n27611) );
  MAO222S U16551 ( .A1(gray_img[489]), .B1(gray_img[488]), .C1(n27451), .O(
        n27452) );
  MAO222S U16552 ( .A1(gray_img[467]), .B1(n26766), .C1(n26765), .O(n26767) );
  MAO222S U16553 ( .A1(n26764), .B1(n26763), .C1(gray_img[466]), .O(n26765) );
  MAO222S U16554 ( .A1(n27570), .B1(gray_img[114]), .C1(n27569), .O(n27571) );
  MAO222S U16555 ( .A1(gray_img[113]), .B1(gray_img[112]), .C1(intadd_122_CI), 
        .O(n27569) );
  MAO222S U16556 ( .A1(n16027), .B1(gray_img[82]), .C1(n16026), .O(n16028) );
  MAO222S U16557 ( .A1(gray_img[81]), .B1(gray_img[80]), .C1(n16025), .O(
        n16026) );
  MAO222 U16558 ( .A1(n26838), .B1(n26836), .C1(n16039), .O(n16040) );
  MAO222 U16559 ( .A1(n23489), .B1(n26845), .C1(n26848), .O(n16039) );
  MAO222S U16560 ( .A1(intadd_171_B_0_), .B1(n23432), .C1(gray_img[129]), .O(
        n23433) );
  OAI12HS U16561 ( .B1(n23906), .B2(n24283), .A1(n23719), .O(n24285) );
  OAI12HS U16562 ( .B1(n23906), .B2(n30456), .A1(n23723), .O(n24319) );
  ND2S U16563 ( .I1(gray_scale_1[5]), .I2(n30444), .O(n19937) );
  AO222S U16564 ( .A1(template_reg[10]), .A2(n17581), .B1(template_reg[2]), 
        .B2(n17579), .C1(n17580), .C2(template_reg[18]), .O(n16096) );
  ND3S U16565 ( .I1(n16094), .I2(n16093), .I3(n16092), .O(n16095) );
  MAO222S U16566 ( .A1(n26548), .B1(gray_img[1554]), .C1(n26547), .O(n26549)
         );
  MAO222S U16567 ( .A1(gray_img[1552]), .B1(gray_img[1553]), .C1(intadd_50_CI), 
        .O(n26547) );
  OR2S U16568 ( .I1(n24679), .I2(n24693), .O(n24684) );
  OR2S U16569 ( .I1(n24680), .I2(n24695), .O(n24683) );
  INV2 U16570 ( .I(n23738), .O(n23736) );
  INV2 U16571 ( .I(n24263), .O(n24328) );
  ND2S U16572 ( .I1(n24835), .I2(n24894), .O(n24807) );
  AO12S U16573 ( .B1(n24198), .B2(n24197), .A1(n24679), .O(n24201) );
  OR2S U16574 ( .I1(n24680), .I2(n15922), .O(n24200) );
  AO12S U16575 ( .B1(n24382), .B2(n24681), .A1(n24346), .O(n24472) );
  OR2S U16576 ( .I1(cnt_cro_3b3[0]), .I2(n24948), .O(n19396) );
  OR2S U16577 ( .I1(n19928), .I2(gray_scale_1[9]), .O(n19932) );
  ND2S U16578 ( .I1(gray_scale_1[7]), .I2(n30450), .O(n19930) );
  INV2 U16579 ( .I(n24429), .O(n24862) );
  MAO222S U16580 ( .A1(n28773), .B1(n28772), .C1(n28771), .O(n28775) );
  MAO222 U16581 ( .A1(n28780), .B1(n28778), .C1(n28770), .O(n28771) );
  MAO222 U16582 ( .A1(n28785), .B1(n28783), .C1(n28769), .O(n28770) );
  MAO222 U16583 ( .A1(n28790), .B1(n28788), .C1(n28768), .O(n28769) );
  MAO222 U16584 ( .A1(gray_img[951]), .B1(n26110), .C1(n26109), .O(n26124) );
  MAO222 U16585 ( .A1(gray_img[950]), .B1(n26108), .C1(n26107), .O(n26109) );
  MAO222 U16586 ( .A1(gray_img[949]), .B1(n26106), .C1(n26105), .O(n26107) );
  MAO222 U16587 ( .A1(gray_img[948]), .B1(n26104), .C1(n26103), .O(n26105) );
  MAO222S U16588 ( .A1(n26132), .B1(n26131), .C1(n26130), .O(n26133) );
  MAO222 U16589 ( .A1(n26135), .B1(n26139), .C1(n26129), .O(n26130) );
  MAO222S U16590 ( .A1(n28255), .B1(n28259), .C1(n26128), .O(n26129) );
  MAO222S U16591 ( .A1(n28221), .B1(n28225), .C1(n26127), .O(n26128) );
  MAO222 U16592 ( .A1(n25969), .B1(gray_img[1911]), .C1(n25968), .O(n25970) );
  MAO222S U16593 ( .A1(n25967), .B1(gray_img[1910]), .C1(n25966), .O(n25968)
         );
  MAO222S U16594 ( .A1(n25965), .B1(gray_img[1909]), .C1(n25964), .O(n25966)
         );
  MAO222 U16595 ( .A1(gray_img[1919]), .B1(n25957), .C1(n25956), .O(n28715) );
  MAO222 U16596 ( .A1(gray_img[1918]), .B1(n25955), .C1(n25954), .O(n25956) );
  MAO222S U16597 ( .A1(n25976), .B1(n25975), .C1(n15969), .O(n25978) );
  AO22S U16598 ( .A1(n25981), .A2(n25983), .B1(n25974), .B2(n15980), .O(n15969) );
  OR2S U16599 ( .I1(n25981), .I2(n25983), .O(n15980) );
  MAO222 U16600 ( .A1(n26057), .B1(n26055), .C1(n15968), .O(n25974) );
  MAO222 U16601 ( .A1(n25848), .B1(gray_img[1895]), .C1(n25847), .O(n25861) );
  MAO222 U16602 ( .A1(n25846), .B1(gray_img[1894]), .C1(n25845), .O(n25847) );
  MAO222 U16603 ( .A1(n25844), .B1(gray_img[1893]), .C1(n25843), .O(n25845) );
  MAO222S U16604 ( .A1(n25842), .B1(gray_img[1892]), .C1(n25841), .O(n25843)
         );
  MAO222 U16605 ( .A1(n25860), .B1(gray_img[1903]), .C1(n25859), .O(n26087) );
  MAO222 U16606 ( .A1(n25858), .B1(gray_img[1902]), .C1(n25857), .O(n25859) );
  MAO222S U16607 ( .A1(n25856), .B1(gray_img[1901]), .C1(n25855), .O(n25857)
         );
  MAO222S U16608 ( .A1(n25854), .B1(gray_img[1900]), .C1(n25853), .O(n25855)
         );
  MAO222S U16609 ( .A1(n25869), .B1(n25868), .C1(n25867), .O(n25871) );
  MAO222 U16610 ( .A1(n25876), .B1(n25874), .C1(n25866), .O(n25867) );
  MAO222 U16611 ( .A1(n25912), .B1(n25910), .C1(n25865), .O(n25866) );
  MAO222 U16612 ( .A1(n25917), .B1(n25915), .C1(n25864), .O(n25865) );
  MAO222 U16613 ( .A1(n24985), .B1(gray_img[815]), .C1(n23219), .O(n23232) );
  MAO222 U16614 ( .A1(n23218), .B1(gray_img[814]), .C1(n23217), .O(n23219) );
  MAO222 U16615 ( .A1(n23216), .B1(gray_img[813]), .C1(n23215), .O(n23217) );
  MAO222 U16616 ( .A1(n23214), .B1(gray_img[812]), .C1(n23213), .O(n23215) );
  MAO222 U16617 ( .A1(n25011), .B1(gray_img[807]), .C1(n23231), .O(n28804) );
  MAO222 U16618 ( .A1(n23230), .B1(gray_img[806]), .C1(n23229), .O(n23231) );
  MAO222S U16619 ( .A1(n23228), .B1(gray_img[805]), .C1(n23227), .O(n23229) );
  MAO222 U16620 ( .A1(gray_img[399]), .B1(n21799), .C1(n18112), .O(n18126) );
  MAO222 U16621 ( .A1(gray_img[398]), .B1(n21225), .C1(n18111), .O(n18112) );
  MAO222 U16622 ( .A1(gray_img[397]), .B1(n18110), .C1(n18109), .O(n18111) );
  MAO222S U16623 ( .A1(n18125), .B1(gray_img[263]), .C1(n18124), .O(n23360) );
  MAO222 U16624 ( .A1(n18123), .B1(gray_img[262]), .C1(n18122), .O(n18124) );
  MAO222 U16625 ( .A1(n18121), .B1(gray_img[261]), .C1(n18120), .O(n18122) );
  MAO222 U16626 ( .A1(n29616), .B1(gray_img[783]), .C1(n29615), .O(n29629) );
  MAO222 U16627 ( .A1(n29614), .B1(gray_img[782]), .C1(n29613), .O(n29615) );
  MAO222 U16628 ( .A1(n29612), .B1(gray_img[781]), .C1(n29611), .O(n29613) );
  MAO222 U16629 ( .A1(n29610), .B1(gray_img[780]), .C1(n29609), .O(n29611) );
  MAO222 U16630 ( .A1(n29628), .B1(gray_img[775]), .C1(n29627), .O(n30100) );
  MAO222S U16631 ( .A1(n29626), .B1(gray_img[774]), .C1(n29625), .O(n29627) );
  MAO222S U16632 ( .A1(n29624), .B1(gray_img[773]), .C1(n29623), .O(n29625) );
  MAO222S U16633 ( .A1(n29637), .B1(n29636), .C1(n29635), .O(n29639) );
  MAO222S U16634 ( .A1(n29644), .B1(n29642), .C1(n29634), .O(n29635) );
  MAO222 U16635 ( .A1(n29975), .B1(n29973), .C1(n29633), .O(n29634) );
  MAO222 U16636 ( .A1(n29980), .B1(n29978), .C1(n29632), .O(n29633) );
  NR2 U16637 ( .I1(n28157), .I2(n28156), .O(n28170) );
  MAO222S U16638 ( .A1(gray_img[702]), .B1(n28153), .C1(n28152), .O(n28155) );
  MAO222 U16639 ( .A1(n28178), .B1(n28177), .C1(n28176), .O(n28179) );
  MAO222 U16640 ( .A1(n28181), .B1(n28185), .C1(n28175), .O(n28176) );
  MAO222 U16641 ( .A1(n28246), .B1(n28254), .C1(n28174), .O(n28175) );
  MAO222S U16642 ( .A1(n28186), .B1(n28190), .C1(n28173), .O(n28174) );
  MAO222 U16643 ( .A1(gray_img[687]), .B1(n28619), .C1(n28618), .O(n28633) );
  MAO222 U16644 ( .A1(gray_img[686]), .B1(n28617), .C1(n28616), .O(n28618) );
  MAO222 U16645 ( .A1(gray_img[685]), .B1(n28615), .C1(n28614), .O(n28616) );
  MAO222S U16646 ( .A1(gray_img[684]), .B1(n28613), .C1(n28612), .O(n28614) );
  MAO222 U16647 ( .A1(n28641), .B1(n28640), .C1(n28639), .O(n28642) );
  MAO222 U16648 ( .A1(n28644), .B1(n28648), .C1(n28638), .O(n28639) );
  MAO222 U16649 ( .A1(n28649), .B1(n28653), .C1(n28637), .O(n28638) );
  MAO222 U16650 ( .A1(n28654), .B1(n28658), .C1(n28636), .O(n28637) );
  MAO222 U16651 ( .A1(n29062), .B1(gray_img[663]), .C1(n29061), .O(n29081) );
  MAO222 U16652 ( .A1(n29060), .B1(gray_img[662]), .C1(n29059), .O(n29061) );
  MAO222S U16653 ( .A1(n29058), .B1(gray_img[661]), .C1(n29057), .O(n29059) );
  MAO222S U16654 ( .A1(n29056), .B1(gray_img[660]), .C1(n29055), .O(n29057) );
  MAO222S U16655 ( .A1(n29089), .B1(n29088), .C1(n29087), .O(n29091) );
  MAO222 U16656 ( .A1(n29096), .B1(n29094), .C1(n29086), .O(n29087) );
  MAO222 U16657 ( .A1(n29319), .B1(n29317), .C1(n29085), .O(n29086) );
  MAO222 U16658 ( .A1(n29329), .B1(n29327), .C1(n29084), .O(n29085) );
  MAO222 U16659 ( .A1(n29917), .B1(gray_img[527]), .C1(n29916), .O(n29930) );
  MAO222 U16660 ( .A1(n29915), .B1(gray_img[526]), .C1(n29914), .O(n29916) );
  MAO222 U16661 ( .A1(n29913), .B1(gray_img[525]), .C1(n29912), .O(n29914) );
  MAO222 U16662 ( .A1(n29929), .B1(gray_img[647]), .C1(n29928), .O(n30002) );
  MAO222S U16663 ( .A1(n29927), .B1(gray_img[646]), .C1(n29926), .O(n29928) );
  MAO222S U16664 ( .A1(n29925), .B1(gray_img[645]), .C1(n29924), .O(n29926) );
  MAO222S U16665 ( .A1(n29923), .B1(gray_img[644]), .C1(n29922), .O(n29924) );
  MAO222S U16666 ( .A1(n29938), .B1(n29937), .C1(n29936), .O(n29940) );
  MAO222S U16667 ( .A1(n29945), .B1(n29943), .C1(n29935), .O(n29936) );
  MAO222S U16668 ( .A1(n29950), .B1(n29948), .C1(n29934), .O(n29935) );
  MAO222S U16669 ( .A1(n29955), .B1(n29953), .C1(n29933), .O(n29934) );
  MAO222 U16670 ( .A1(n27863), .B1(gray_img[151]), .C1(n27862), .O(n30078) );
  MAO222 U16671 ( .A1(n27861), .B1(gray_img[150]), .C1(n27860), .O(n27862) );
  MAO222 U16672 ( .A1(n27859), .B1(gray_img[149]), .C1(n27858), .O(n27860) );
  MAO222 U16673 ( .A1(n27876), .B1(gray_img[31]), .C1(n27875), .O(n27877) );
  MAO222 U16674 ( .A1(n27874), .B1(gray_img[30]), .C1(n27873), .O(n27875) );
  MAO222 U16675 ( .A1(n27872), .B1(gray_img[29]), .C1(n27871), .O(n27873) );
  MAO222 U16676 ( .A1(n27870), .B1(gray_img[28]), .C1(n27869), .O(n27871) );
  MAO222 U16677 ( .A1(n26501), .B1(gray_img[447]), .C1(n26500), .O(n26514) );
  MAO222 U16678 ( .A1(n26499), .B1(gray_img[446]), .C1(n26498), .O(n26500) );
  MAO222 U16679 ( .A1(n26497), .B1(gray_img[445]), .C1(n26496), .O(n26498) );
  MAO222 U16680 ( .A1(n26513), .B1(gray_img[439]), .C1(n26512), .O(n27842) );
  MAO222 U16681 ( .A1(n26511), .B1(gray_img[438]), .C1(n26510), .O(n26512) );
  MAO222S U16682 ( .A1(n26509), .B1(gray_img[437]), .C1(n26508), .O(n26510) );
  MAO222S U16683 ( .A1(n26521), .B1(n26520), .C1(n26519), .O(n26523) );
  MAO222 U16684 ( .A1(n26528), .B1(n26526), .C1(n26518), .O(n26519) );
  MAO222 U16685 ( .A1(n27798), .B1(n27796), .C1(n26517), .O(n26518) );
  MAO222S U16686 ( .A1(n27803), .B1(n27801), .C1(n15978), .O(n26517) );
  MAO222 U16687 ( .A1(n27287), .B1(gray_img[431]), .C1(n27286), .O(n30067) );
  MAO222 U16688 ( .A1(n27285), .B1(gray_img[430]), .C1(n27284), .O(n27286) );
  MAO222 U16689 ( .A1(n27275), .B1(gray_img[423]), .C1(n27274), .O(n27288) );
  MAO222 U16690 ( .A1(n27273), .B1(gray_img[422]), .C1(n27272), .O(n27274) );
  MAO222 U16691 ( .A1(n27271), .B1(gray_img[421]), .C1(n27270), .O(n27272) );
  MAO222S U16692 ( .A1(n27296), .B1(n27295), .C1(n27294), .O(n27298) );
  MAO222S U16693 ( .A1(n27303), .B1(n27301), .C1(n27293), .O(n27294) );
  MAO222S U16694 ( .A1(n27308), .B1(n27306), .C1(n27292), .O(n27293) );
  MAO222 U16695 ( .A1(n27313), .B1(n27311), .C1(n27291), .O(n27292) );
  MAO222S U16696 ( .A1(n27743), .B1(n27742), .C1(n27741), .O(n27745) );
  MAO222 U16697 ( .A1(n27761), .B1(n27759), .C1(n27738), .O(n27739) );
  MAO222 U16698 ( .A1(n26955), .B1(gray_img[39]), .C1(n26954), .O(n26969) );
  MAO222 U16699 ( .A1(n26953), .B1(gray_img[38]), .C1(n26952), .O(n26954) );
  MAO222S U16700 ( .A1(n26951), .B1(gray_img[37]), .C1(n26950), .O(n26952) );
  MAO222 U16701 ( .A1(n26968), .B1(gray_img[175]), .C1(n26967), .O(n27363) );
  MAO222S U16702 ( .A1(n26966), .B1(gray_img[174]), .C1(n26965), .O(n26967) );
  MAO222S U16703 ( .A1(n26964), .B1(gray_img[173]), .C1(n26963), .O(n26965) );
  MAO222 U16704 ( .A1(n26977), .B1(n26976), .C1(n26975), .O(n26979) );
  MAO222 U16705 ( .A1(n26984), .B1(n26982), .C1(n26974), .O(n26975) );
  MAO222 U16706 ( .A1(n27334), .B1(n27332), .C1(n26973), .O(n26974) );
  MAO222 U16707 ( .A1(n27339), .B1(n27337), .C1(n26972), .O(n26973) );
  MAO222 U16708 ( .A1(n25001), .B1(gray_img[1871]), .C1(n23572), .O(n23582) );
  MAO222 U16709 ( .A1(n23571), .B1(gray_img[1870]), .C1(n23570), .O(n23572) );
  MAO222 U16710 ( .A1(n23569), .B1(gray_img[1869]), .C1(n23568), .O(n23570) );
  MAO222 U16711 ( .A1(n23567), .B1(gray_img[1868]), .C1(n23566), .O(n23568) );
  MAO222 U16712 ( .A1(gray_img[1863]), .B1(n23560), .C1(n23559), .O(n23573) );
  MAO222 U16713 ( .A1(gray_img[1862]), .B1(n23558), .C1(n23557), .O(n23559) );
  MAO222 U16714 ( .A1(gray_img[1861]), .B1(n23556), .C1(n23555), .O(n23557) );
  MAO222S U16715 ( .A1(gray_img[1860]), .B1(n23554), .C1(n23553), .O(n23555)
         );
  MAO222S U16716 ( .A1(n29298), .B1(gray_img[791]), .C1(n29297), .O(n30029) );
  MAO222 U16717 ( .A1(n29296), .B1(gray_img[790]), .C1(n29295), .O(n29297) );
  MAO222 U16718 ( .A1(n29286), .B1(gray_img[799]), .C1(n29285), .O(n29299) );
  MAO222 U16719 ( .A1(n29284), .B1(gray_img[798]), .C1(n29283), .O(n29285) );
  MAO222S U16720 ( .A1(n29282), .B1(gray_img[797]), .C1(n29281), .O(n29283) );
  MAO222 U16721 ( .A1(n29307), .B1(n29306), .C1(n29305), .O(n29309) );
  MAO222S U16722 ( .A1(n29314), .B1(n29312), .C1(n29304), .O(n29305) );
  MAO222S U16723 ( .A1(n29324), .B1(n29322), .C1(n29303), .O(n29304) );
  MAO222 U16724 ( .A1(n29363), .B1(n29361), .C1(n29302), .O(n29303) );
  MAO222 U16725 ( .A1(n23138), .B1(gray_img[1855]), .C1(n23137), .O(n23151) );
  MAO222 U16726 ( .A1(n23136), .B1(gray_img[1854]), .C1(n23135), .O(n23137) );
  MAO222S U16727 ( .A1(n23134), .B1(gray_img[1853]), .C1(n23133), .O(n23135)
         );
  MAO222 U16728 ( .A1(n23150), .B1(gray_img[1847]), .C1(n23149), .O(n23162) );
  MAO222 U16729 ( .A1(n23148), .B1(gray_img[1846]), .C1(n23147), .O(n23149) );
  MAO222 U16730 ( .A1(n23146), .B1(gray_img[1845]), .C1(n23145), .O(n23147) );
  MAO222 U16731 ( .A1(gray_img[1831]), .B1(n26668), .C1(n26667), .O(n26682) );
  MAO222 U16732 ( .A1(gray_img[1830]), .B1(n26666), .C1(n26665), .O(n26667) );
  MAO222 U16733 ( .A1(gray_img[1829]), .B1(n26664), .C1(n26663), .O(n26665) );
  MAO222 U16734 ( .A1(gray_img[1828]), .B1(n26662), .C1(n26661), .O(n26663) );
  MAO222S U16735 ( .A1(n26690), .B1(n26689), .C1(n26688), .O(n26691) );
  MAO222 U16736 ( .A1(n26693), .B1(n26697), .C1(n26687), .O(n26688) );
  MAO222 U16737 ( .A1(n29162), .B1(n29166), .C1(n26686), .O(n26687) );
  MAO222 U16738 ( .A1(n29167), .B1(n29171), .C1(n26685), .O(n26686) );
  MAO222 U16739 ( .A1(n29516), .B1(gray_img[1823]), .C1(n29515), .O(n29517) );
  MAO222 U16740 ( .A1(n29514), .B1(gray_img[1822]), .C1(n29513), .O(n29515) );
  MAO222 U16741 ( .A1(n29512), .B1(gray_img[1821]), .C1(n29511), .O(n29513) );
  MAO222S U16742 ( .A1(n29504), .B1(gray_img[1815]), .C1(n29503), .O(n29594)
         );
  MAO222 U16743 ( .A1(n29502), .B1(gray_img[1814]), .C1(n29501), .O(n29503) );
  MAO222S U16744 ( .A1(n29523), .B1(n29522), .C1(n15954), .O(n29525) );
  AO22S U16745 ( .A1(n29528), .A2(n29530), .B1(n29521), .B2(n15972), .O(n15954) );
  OR2S U16746 ( .I1(n29528), .I2(n29530), .O(n15972) );
  MAO222 U16747 ( .A1(n29560), .B1(n29558), .C1(n15953), .O(n29521) );
  MAO222 U16748 ( .A1(n29399), .B1(gray_img[1927]), .C1(n29398), .O(n30089) );
  MAO222 U16749 ( .A1(n29397), .B1(gray_img[1926]), .C1(n29396), .O(n29398) );
  MAO222S U16750 ( .A1(n29395), .B1(gray_img[1925]), .C1(n29394), .O(n29396)
         );
  MAO222S U16751 ( .A1(n29393), .B1(gray_img[1924]), .C1(n29392), .O(n29394)
         );
  MOAI1S U16752 ( .A1(gray_img[1806]), .A2(n29410), .B1(n29409), .B2(
        gray_img[1934]), .O(n29413) );
  ND2S U16753 ( .I1(n29410), .I2(gray_img[1806]), .O(n29409) );
  MAO222 U16754 ( .A1(n29423), .B1(n29422), .C1(n29421), .O(n29424) );
  MAO222S U16755 ( .A1(n29426), .B1(n29431), .C1(n29420), .O(n29421) );
  MAO222 U16756 ( .A1(n29461), .B1(n29459), .C1(n29419), .O(n29420) );
  MAO222 U16757 ( .A1(n29466), .B1(n29464), .C1(n29418), .O(n29419) );
  MAO222 U16758 ( .A1(n25995), .B1(gray_img[1663]), .C1(n25994), .O(n26009) );
  MAO222 U16759 ( .A1(n25993), .B1(gray_img[1662]), .C1(n25992), .O(n25994) );
  MAO222 U16760 ( .A1(n25991), .B1(gray_img[1661]), .C1(n25990), .O(n25992) );
  MAO222 U16761 ( .A1(n26008), .B1(gray_img[1655]), .C1(n26007), .O(n26045) );
  MAO222S U16762 ( .A1(n26006), .B1(gray_img[1654]), .C1(n26005), .O(n26007)
         );
  MAO222S U16763 ( .A1(n26017), .B1(n26016), .C1(n26015), .O(n26019) );
  MAO222 U16764 ( .A1(n26024), .B1(n26022), .C1(n26014), .O(n26015) );
  MAO222 U16765 ( .A1(n26029), .B1(n26027), .C1(n26013), .O(n26014) );
  MAO222 U16766 ( .A1(n26034), .B1(n26032), .C1(n26012), .O(n26013) );
  MAO222S U16767 ( .A1(n25804), .B1(gray_img[1767]), .C1(n25803), .O(n25900)
         );
  MAO222 U16768 ( .A1(n25802), .B1(gray_img[1766]), .C1(n25801), .O(n25803) );
  MAO222 U16769 ( .A1(n25800), .B1(gray_img[1765]), .C1(n25799), .O(n25801) );
  MAO222 U16770 ( .A1(n25792), .B1(gray_img[1775]), .C1(n25791), .O(n25805) );
  MAO222S U16771 ( .A1(n25790), .B1(gray_img[1774]), .C1(n25789), .O(n25791)
         );
  MAO222S U16772 ( .A1(n25788), .B1(gray_img[1773]), .C1(n25787), .O(n25789)
         );
  MAO222S U16773 ( .A1(n25786), .B1(gray_img[1772]), .C1(n25785), .O(n25787)
         );
  MAO222S U16774 ( .A1(n25813), .B1(n25812), .C1(n25811), .O(n25815) );
  MAO222S U16775 ( .A1(n25820), .B1(n25818), .C1(n25810), .O(n25811) );
  MAO222 U16776 ( .A1(n25881), .B1(n25879), .C1(n25809), .O(n25810) );
  MAO222 U16777 ( .A1(n25886), .B1(n25884), .C1(n25808), .O(n25809) );
  MAO222 U16778 ( .A1(gray_img[1751]), .B1(n25524), .C1(n25523), .O(n25538) );
  MAO222S U16779 ( .A1(gray_img[1750]), .B1(n25522), .C1(n25521), .O(n25523)
         );
  MAO222 U16780 ( .A1(gray_img[1749]), .B1(n25520), .C1(n25519), .O(n25521) );
  MAO222 U16781 ( .A1(gray_img[1748]), .B1(n25518), .C1(n25517), .O(n25519) );
  MAO222 U16782 ( .A1(n25546), .B1(n25545), .C1(n25544), .O(n25547) );
  MAO222S U16783 ( .A1(n25549), .B1(n25553), .C1(n25543), .O(n25544) );
  MAO222S U16784 ( .A1(n25554), .B1(n25558), .C1(n25542), .O(n25543) );
  MAO222S U16785 ( .A1(n25559), .B1(n25563), .C1(n25541), .O(n25542) );
  MAO222 U16786 ( .A1(n25678), .B1(gray_img[1735]), .C1(n25677), .O(n25741) );
  MAO222 U16787 ( .A1(n25676), .B1(gray_img[1734]), .C1(n25675), .O(n25677) );
  MAO222 U16788 ( .A1(n25674), .B1(gray_img[1733]), .C1(n25673), .O(n25675) );
  MAO222 U16789 ( .A1(n25666), .B1(gray_img[1743]), .C1(n25665), .O(n25679) );
  MAO222 U16790 ( .A1(n25664), .B1(gray_img[1742]), .C1(n25663), .O(n25665) );
  MAO222S U16791 ( .A1(n25662), .B1(gray_img[1741]), .C1(n25661), .O(n25663)
         );
  MAO222S U16792 ( .A1(n25660), .B1(gray_img[1740]), .C1(n25659), .O(n25661)
         );
  MAO222S U16793 ( .A1(n25687), .B1(n25686), .C1(n25685), .O(n25689) );
  MAO222S U16794 ( .A1(n25694), .B1(n25692), .C1(n25684), .O(n25685) );
  MAO222 U16795 ( .A1(n25699), .B1(n25697), .C1(n25683), .O(n25684) );
  MAO222 U16796 ( .A1(n25704), .B1(n25702), .C1(n25682), .O(n25683) );
  MAO222 U16797 ( .A1(n29209), .B1(gray_img[1599]), .C1(n29208), .O(n29258) );
  MAO222 U16798 ( .A1(n29207), .B1(gray_img[1598]), .C1(n29206), .O(n29208) );
  MAO222 U16799 ( .A1(n29205), .B1(gray_img[1597]), .C1(n29204), .O(n29206) );
  MAO222 U16800 ( .A1(n29221), .B1(gray_img[1591]), .C1(n29220), .O(n29222) );
  MAO222 U16801 ( .A1(n29219), .B1(gray_img[1590]), .C1(n29218), .O(n29220) );
  MAO222 U16802 ( .A1(n29217), .B1(gray_img[1589]), .C1(n29216), .O(n29218) );
  MAO222S U16803 ( .A1(n29230), .B1(n29229), .C1(n29228), .O(n29231) );
  MAO222 U16804 ( .A1(n29233), .B1(n29237), .C1(n29227), .O(n29228) );
  MAO222 U16805 ( .A1(n29242), .B1(n29240), .C1(n29226), .O(n29227) );
  MAO222 U16806 ( .A1(n29247), .B1(n29245), .C1(n29225), .O(n29226) );
  MAO222S U16807 ( .A1(n29108), .B1(gray_img[1583]), .C1(n29107), .O(n29121)
         );
  MAO222 U16808 ( .A1(n29106), .B1(gray_img[1582]), .C1(n29105), .O(n29107) );
  MAO222 U16809 ( .A1(n29104), .B1(gray_img[1581]), .C1(n29103), .O(n29105) );
  MAO222S U16810 ( .A1(n29120), .B1(gray_img[1575]), .C1(n29119), .O(n29183)
         );
  MAO222 U16811 ( .A1(n29118), .B1(gray_img[1574]), .C1(n29117), .O(n29119) );
  MAO222S U16812 ( .A1(n29129), .B1(n29128), .C1(n29127), .O(n29131) );
  MAO222 U16813 ( .A1(n29136), .B1(n29134), .C1(n29126), .O(n29127) );
  MAO222S U16814 ( .A1(n29141), .B1(n29139), .C1(n29125), .O(n29126) );
  MAO222 U16815 ( .A1(n29146), .B1(n29144), .C1(n29124), .O(n29125) );
  OAI12HS U16816 ( .B1(gray_img[1695]), .B2(n26546), .A1(n26545), .O(n26559)
         );
  MAO222 U16817 ( .A1(n26567), .B1(n26566), .C1(n26565), .O(n26568) );
  MAO222 U16818 ( .A1(n26570), .B1(n26574), .C1(n26564), .O(n26565) );
  MAO222 U16819 ( .A1(n29531), .B1(n29535), .C1(n26563), .O(n26564) );
  MAO222 U16820 ( .A1(n29536), .B1(n29540), .C1(n26562), .O(n26563) );
  MAO222 U16821 ( .A1(n26600), .B1(gray_img[1671]), .C1(n26599), .O(n29478) );
  MAO222S U16822 ( .A1(n26598), .B1(gray_img[1670]), .C1(n26597), .O(n26599)
         );
  MAO222 U16823 ( .A1(n26596), .B1(gray_img[1669]), .C1(n26595), .O(n26597) );
  MAO222 U16824 ( .A1(n26594), .B1(gray_img[1668]), .C1(n26593), .O(n26595) );
  MAO222 U16825 ( .A1(n26587), .B1(gray_img[1551]), .C1(n26586), .O(n26601) );
  MAO222 U16826 ( .A1(n26585), .B1(gray_img[1550]), .C1(n26584), .O(n26586) );
  MAO222S U16827 ( .A1(n26583), .B1(gray_img[1549]), .C1(n26582), .O(n26584)
         );
  MAO222 U16828 ( .A1(n26609), .B1(n26608), .C1(n26607), .O(n26611) );
  MAO222 U16829 ( .A1(n26616), .B1(n26614), .C1(n26606), .O(n26607) );
  MAO222 U16830 ( .A1(n29436), .B1(n29434), .C1(n26605), .O(n26606) );
  MAO222 U16831 ( .A1(n29441), .B1(n29439), .C1(n26604), .O(n26605) );
  MAO222 U16832 ( .A1(n27904), .B1(gray_img[1407]), .C1(n27903), .O(n27918) );
  MAO222 U16833 ( .A1(n27902), .B1(gray_img[1406]), .C1(n27901), .O(n27903) );
  MAO222 U16834 ( .A1(n27984), .B1(gray_img[1391]), .C1(n27983), .O(n28003) );
  MAO222 U16835 ( .A1(n27982), .B1(gray_img[1390]), .C1(n27981), .O(n27983) );
  MAO222 U16836 ( .A1(n27980), .B1(gray_img[1389]), .C1(n27979), .O(n27981) );
  ND3S U16837 ( .I1(n28000), .I2(n27999), .I3(n27998), .O(n28001) );
  MAO222S U16838 ( .A1(n28011), .B1(n28010), .C1(n28009), .O(n28013) );
  MAO222 U16839 ( .A1(n28018), .B1(n28016), .C1(n28008), .O(n28009) );
  MAO222 U16840 ( .A1(n28105), .B1(n28103), .C1(n28007), .O(n28008) );
  MAO222S U16841 ( .A1(n28110), .B1(n28108), .C1(n28006), .O(n28007) );
  MAO222 U16842 ( .A1(n28384), .B1(gray_img[1495]), .C1(n28383), .O(n28598) );
  MAO222 U16843 ( .A1(n28382), .B1(gray_img[1494]), .C1(n28381), .O(n28383) );
  MAO222 U16844 ( .A1(n28372), .B1(gray_img[1503]), .C1(n28371), .O(n28385) );
  MAO222 U16845 ( .A1(n28370), .B1(gray_img[1502]), .C1(n28369), .O(n28371) );
  MAO222 U16846 ( .A1(n28368), .B1(gray_img[1501]), .C1(n28367), .O(n28369) );
  MAO222S U16847 ( .A1(n28393), .B1(n28392), .C1(n28391), .O(n28395) );
  MAO222S U16848 ( .A1(n28400), .B1(n28398), .C1(n28390), .O(n28391) );
  MAO222 U16849 ( .A1(n28436), .B1(n28434), .C1(n28389), .O(n28390) );
  MAO222 U16850 ( .A1(n28441), .B1(n28439), .C1(n28388), .O(n28389) );
  NR2 U16851 ( .I1(n23514), .I2(n23513), .O(n23530) );
  MAO222 U16852 ( .A1(gray_img[1350]), .B1(n23510), .C1(n23509), .O(n23512) );
  MAO222 U16853 ( .A1(n21934), .B1(gray_img[1343]), .C1(n18065), .O(n29341) );
  MAO222 U16854 ( .A1(n18064), .B1(gray_img[1342]), .C1(n18063), .O(n18065) );
  MAO222 U16855 ( .A1(n18062), .B1(gray_img[1341]), .C1(n18061), .O(n18063) );
  MOAI1S U16856 ( .A1(n18083), .A2(n18082), .B1(gray_img[1335]), .B2(n18081), 
        .O(n18084) );
  MAO222S U16857 ( .A1(n25311), .B1(n25312), .C1(n18090), .O(n18091) );
  MAO222 U16858 ( .A1(n18093), .B1(n18101), .C1(n18089), .O(n18090) );
  MAO222S U16859 ( .A1(n28899), .B1(n28897), .C1(n18088), .O(n18089) );
  MAO222 U16860 ( .A1(n23202), .B1(n23205), .C1(n18087), .O(n18088) );
  MAO222 U16861 ( .A1(n28974), .B1(gray_img[1327]), .C1(n28973), .O(n28975) );
  MAO222 U16862 ( .A1(n28972), .B1(gray_img[1326]), .C1(n28971), .O(n28973) );
  MAO222S U16863 ( .A1(n28970), .B1(gray_img[1325]), .C1(n28969), .O(n28971)
         );
  MAO222 U16864 ( .A1(n28962), .B1(gray_img[1319]), .C1(n28961), .O(n29009) );
  MAO222 U16865 ( .A1(n28960), .B1(gray_img[1318]), .C1(n28959), .O(n28961) );
  MAO222 U16866 ( .A1(n28958), .B1(gray_img[1317]), .C1(n28957), .O(n28959) );
  MAO222S U16867 ( .A1(n28981), .B1(n28980), .C1(n15973), .O(n28983) );
  AO22S U16868 ( .A1(n28986), .A2(n28988), .B1(n28979), .B2(n15967), .O(n15973) );
  OR2S U16869 ( .I1(n28986), .I2(n28988), .O(n15967) );
  MAO222 U16870 ( .A1(n28993), .B1(n28991), .C1(n15966), .O(n28979) );
  MAO222 U16871 ( .A1(n29759), .B1(gray_img[1431]), .C1(n29758), .O(n29773) );
  MAO222S U16872 ( .A1(n29757), .B1(gray_img[1430]), .C1(n29756), .O(n29758)
         );
  MAO222S U16873 ( .A1(n29755), .B1(gray_img[1429]), .C1(n29754), .O(n29756)
         );
  MAO222S U16874 ( .A1(n29753), .B1(gray_img[1428]), .C1(n29752), .O(n29754)
         );
  MAO222 U16875 ( .A1(n29772), .B1(gray_img[1439]), .C1(n29771), .O(n29895) );
  MAO222 U16876 ( .A1(n29770), .B1(gray_img[1438]), .C1(n29769), .O(n29771) );
  MAO222S U16877 ( .A1(n29768), .B1(gray_img[1437]), .C1(n29767), .O(n29769)
         );
  MAO222 U16878 ( .A1(n29781), .B1(n29780), .C1(n29779), .O(n29783) );
  MAO222 U16879 ( .A1(n29788), .B1(n29786), .C1(n29778), .O(n29779) );
  MAO222S U16880 ( .A1(n29863), .B1(n29861), .C1(n29777), .O(n29778) );
  MAO222 U16881 ( .A1(n29868), .B1(n29866), .C1(n29776), .O(n29777) );
  MAO222 U16882 ( .A1(n29656), .B1(gray_img[1287]), .C1(n29655), .O(n29669) );
  MAO222 U16883 ( .A1(n29654), .B1(gray_img[1286]), .C1(n29653), .O(n29655) );
  MAO222 U16884 ( .A1(n29652), .B1(gray_img[1285]), .C1(n29651), .O(n29653) );
  MAO222 U16885 ( .A1(n29677), .B1(n29676), .C1(n29675), .O(n29678) );
  MAO222 U16886 ( .A1(n29681), .B1(n29685), .C1(n29674), .O(n29675) );
  MAO222 U16887 ( .A1(n29686), .B1(n29690), .C1(n29673), .O(n29674) );
  MAO222 U16888 ( .A1(n29691), .B1(n29695), .C1(n29672), .O(n29673) );
  MAO222 U16889 ( .A1(n23311), .B1(gray_img[1271]), .C1(n23310), .O(n23324) );
  MAO222 U16890 ( .A1(n23309), .B1(gray_img[1270]), .C1(n23308), .O(n23310) );
  MAO222 U16891 ( .A1(n23307), .B1(gray_img[1269]), .C1(n23306), .O(n23308) );
  MAO222 U16892 ( .A1(n23323), .B1(gray_img[1151]), .C1(n23322), .O(n23490) );
  MAO222 U16893 ( .A1(n23321), .B1(gray_img[1150]), .C1(n23320), .O(n23322) );
  MAO222 U16894 ( .A1(n23319), .B1(gray_img[1149]), .C1(n23318), .O(n23320) );
  MAO222 U16895 ( .A1(n28055), .B1(gray_img[1263]), .C1(n28054), .O(n28056) );
  MAO222 U16896 ( .A1(n28053), .B1(gray_img[1262]), .C1(n28052), .O(n28054) );
  MAO222S U16897 ( .A1(n28051), .B1(gray_img[1261]), .C1(n28050), .O(n28052)
         );
  MAO222S U16898 ( .A1(n28049), .B1(gray_img[1260]), .C1(n28048), .O(n28050)
         );
  MAO222S U16899 ( .A1(n28043), .B1(gray_img[1127]), .C1(n28042), .O(n28093)
         );
  MAO222S U16900 ( .A1(n28041), .B1(gray_img[1126]), .C1(n28040), .O(n28042)
         );
  MAO222 U16901 ( .A1(n28039), .B1(gray_img[1125]), .C1(n28038), .O(n28040) );
  MAO222 U16902 ( .A1(n28037), .B1(gray_img[1124]), .C1(n28036), .O(n28038) );
  MAO222S U16903 ( .A1(n28062), .B1(n28061), .C1(n15956), .O(n28064) );
  AO22S U16904 ( .A1(n28067), .A2(n28069), .B1(n28060), .B2(n15964), .O(n15956) );
  OR2S U16905 ( .I1(n28067), .I2(n28069), .O(n15964) );
  MAO222 U16906 ( .A1(n28074), .B1(n28072), .C1(n15955), .O(n28060) );
  MAO222 U16907 ( .A1(n28301), .B1(gray_img[1119]), .C1(n28300), .O(n28315) );
  MAO222S U16908 ( .A1(n28299), .B1(gray_img[1118]), .C1(n28298), .O(n28300)
         );
  MAO222 U16909 ( .A1(n28297), .B1(gray_img[1117]), .C1(n28296), .O(n28298) );
  MAO222 U16910 ( .A1(n28314), .B1(gray_img[1239]), .C1(n28313), .O(n28424) );
  MAO222 U16911 ( .A1(n28312), .B1(gray_img[1238]), .C1(n28311), .O(n28313) );
  MAO222S U16912 ( .A1(n28323), .B1(n28322), .C1(n28321), .O(n28325) );
  MAO222S U16913 ( .A1(n28330), .B1(n28328), .C1(n28320), .O(n28321) );
  MAO222 U16914 ( .A1(n28405), .B1(n28403), .C1(n28319), .O(n28320) );
  MAO222 U16915 ( .A1(n28410), .B1(n28408), .C1(n28318), .O(n28319) );
  MAO222 U16916 ( .A1(gray_img[1103]), .B1(n28494), .C1(n28493), .O(n28507) );
  MAO222 U16917 ( .A1(gray_img[1102]), .B1(n28492), .C1(n28491), .O(n28493) );
  MAO222 U16918 ( .A1(n28515), .B1(n28514), .C1(n28513), .O(n28516) );
  MAO222 U16919 ( .A1(n28518), .B1(n28522), .C1(n28512), .O(n28513) );
  MAO222 U16920 ( .A1(n28561), .B1(n28565), .C1(n28511), .O(n28512) );
  MAO222 U16921 ( .A1(n28566), .B1(n28570), .C1(n28510), .O(n28511) );
  MAO222 U16922 ( .A1(n28865), .B1(gray_img[1087]), .C1(n28864), .O(n28879) );
  MAO222 U16923 ( .A1(n28863), .B1(gray_img[1086]), .C1(n28862), .O(n28864) );
  MAO222S U16924 ( .A1(n28861), .B1(gray_img[1085]), .C1(n28860), .O(n28862)
         );
  MAO222S U16925 ( .A1(n28878), .B1(gray_img[1079]), .C1(n28877), .O(n28935)
         );
  MAO222 U16926 ( .A1(n28876), .B1(gray_img[1078]), .C1(n28875), .O(n28877) );
  MAO222 U16927 ( .A1(n28874), .B1(gray_img[1077]), .C1(n28873), .O(n28875) );
  MAO222S U16928 ( .A1(n28887), .B1(n28886), .C1(n28885), .O(n28889) );
  MAO222S U16929 ( .A1(n28894), .B1(n28892), .C1(n28884), .O(n28885) );
  MAO222 U16930 ( .A1(n28904), .B1(n28902), .C1(n28883), .O(n28884) );
  MAO222 U16931 ( .A1(n28924), .B1(n28922), .C1(n28882), .O(n28883) );
  MAO222 U16932 ( .A1(n23020), .B1(gray_img[1063]), .C1(n23019), .O(n23033) );
  MAO222 U16933 ( .A1(n23018), .B1(gray_img[1062]), .C1(n23017), .O(n23019) );
  MAO222 U16934 ( .A1(n23016), .B1(gray_img[1061]), .C1(n23015), .O(n23017) );
  MAO222S U16935 ( .A1(n23014), .B1(gray_img[1060]), .C1(n23013), .O(n23015)
         );
  MAO222 U16936 ( .A1(n23032), .B1(gray_img[1071]), .C1(n23031), .O(n29041) );
  MAO222 U16937 ( .A1(n23030), .B1(gray_img[1070]), .C1(n23029), .O(n23031) );
  MAO222S U16938 ( .A1(n23028), .B1(gray_img[1069]), .C1(n23027), .O(n23029)
         );
  MAO222 U16939 ( .A1(n23041), .B1(n23040), .C1(n23039), .O(n23042) );
  MAO222S U16940 ( .A1(n26140), .B1(n26144), .C1(n23038), .O(n23039) );
  MAO222S U16941 ( .A1(n29017), .B1(n29021), .C1(n23037), .O(n23038) );
  MAO222 U16942 ( .A1(n29022), .B1(n29026), .C1(n23036), .O(n23037) );
  MAO222 U16943 ( .A1(n29799), .B1(gray_img[1055]), .C1(n29798), .O(n29812) );
  MAO222 U16944 ( .A1(n29797), .B1(gray_img[1054]), .C1(n29796), .O(n29798) );
  MAO222 U16945 ( .A1(n29795), .B1(gray_img[1053]), .C1(n29794), .O(n29796) );
  MAO222 U16946 ( .A1(n29811), .B1(gray_img[1047]), .C1(n29810), .O(n29853) );
  MAO222 U16947 ( .A1(n29809), .B1(gray_img[1046]), .C1(n29808), .O(n29810) );
  MAO222 U16948 ( .A1(n29807), .B1(gray_img[1045]), .C1(n29806), .O(n29808) );
  MAO222 U16949 ( .A1(n29820), .B1(n29819), .C1(n29818), .O(n29821) );
  MAO222 U16950 ( .A1(n29823), .B1(n29828), .C1(n29817), .O(n29818) );
  MAO222 U16951 ( .A1(n29829), .B1(n29834), .C1(n29816), .O(n29817) );
  MAO222 U16952 ( .A1(n29835), .B1(n29840), .C1(n29815), .O(n29816) );
  MAO222 U16953 ( .A1(n26627), .B1(gray_img[1167]), .C1(n26626), .O(n26640) );
  MAO222 U16954 ( .A1(n26625), .B1(gray_img[1166]), .C1(n26624), .O(n26626) );
  MAO222 U16955 ( .A1(n26623), .B1(gray_img[1165]), .C1(n26622), .O(n26624) );
  MAO222S U16956 ( .A1(n26621), .B1(gray_img[1164]), .C1(n26620), .O(n26622)
         );
  MAO222 U16957 ( .A1(n26648), .B1(n26647), .C1(n26646), .O(n26649) );
  MAO222 U16958 ( .A1(n26651), .B1(n26655), .C1(n26645), .O(n26646) );
  MAO222 U16959 ( .A1(n29711), .B1(n29715), .C1(n26644), .O(n26645) );
  MAO222 U16960 ( .A1(n29716), .B1(n29720), .C1(n26643), .O(n26644) );
  MAO222 U16961 ( .A1(n26387), .B1(gray_img[1015]), .C1(n26386), .O(n26401) );
  MAO222 U16962 ( .A1(n26385), .B1(gray_img[1014]), .C1(n26384), .O(n26386) );
  MAO222 U16963 ( .A1(n26383), .B1(gray_img[1013]), .C1(n26382), .O(n26384) );
  MAO222S U16964 ( .A1(n26381), .B1(gray_img[1012]), .C1(n26380), .O(n26382)
         );
  MAO222 U16965 ( .A1(n26400), .B1(gray_img[1023]), .C1(n26399), .O(n26437) );
  MAO222S U16966 ( .A1(n26398), .B1(gray_img[1022]), .C1(n26397), .O(n26399)
         );
  MAO222S U16967 ( .A1(n26409), .B1(n26408), .C1(n26407), .O(n26411) );
  MAO222 U16968 ( .A1(n26416), .B1(n26414), .C1(n26406), .O(n26407) );
  MAO222 U16969 ( .A1(n26421), .B1(n26419), .C1(n26405), .O(n26406) );
  MAO222 U16970 ( .A1(n26426), .B1(n26424), .C1(n26404), .O(n26405) );
  MAO222 U16971 ( .A1(n26255), .B1(gray_img[871]), .C1(n26254), .O(n27831) );
  MAO222 U16972 ( .A1(n26253), .B1(gray_img[870]), .C1(n26252), .O(n26254) );
  MAO222 U16973 ( .A1(n26251), .B1(gray_img[869]), .C1(n26250), .O(n26252) );
  MAO222S U16974 ( .A1(n26264), .B1(n26263), .C1(n26262), .O(n26266) );
  MAO222S U16975 ( .A1(n26271), .B1(n26269), .C1(n26261), .O(n26262) );
  MAO222 U16976 ( .A1(n26276), .B1(n26274), .C1(n26260), .O(n26261) );
  MAO222S U16977 ( .A1(n26281), .B1(n26279), .C1(n26259), .O(n26260) );
  MAO222 U16978 ( .A1(n23066), .B1(gray_img[983]), .C1(n23065), .O(n23079) );
  MAO222 U16979 ( .A1(n23064), .B1(gray_img[982]), .C1(n23063), .O(n23065) );
  MAO222 U16980 ( .A1(n23062), .B1(gray_img[981]), .C1(n23061), .O(n23063) );
  MAO222 U16981 ( .A1(n23078), .B1(gray_img[991]), .C1(n23077), .O(n23088) );
  MAO222 U16982 ( .A1(n23076), .B1(gray_img[990]), .C1(n23075), .O(n23077) );
  MAO222 U16983 ( .A1(n23074), .B1(gray_img[989]), .C1(n23073), .O(n23075) );
  MAO222 U16984 ( .A1(n23072), .B1(gray_img[988]), .C1(n23071), .O(n23073) );
  MAO222S U16985 ( .A1(n25148), .B1(n25149), .C1(n23085), .O(n23086) );
  MAO222 U16986 ( .A1(n23115), .B1(n23119), .C1(n23084), .O(n23085) );
  MAO222 U16987 ( .A1(n23110), .B1(n23114), .C1(n23083), .O(n23084) );
  MAO222 U16988 ( .A1(n23105), .B1(n23109), .C1(n23082), .O(n23083) );
  MAO222 U16989 ( .A1(n23002), .B1(n23001), .C1(n23000), .O(n23004) );
  ND2S U16990 ( .I1(n22997), .I2(n22996), .O(n22998) );
  MAO222S U16991 ( .A1(n22995), .B1(n23008), .C1(n23005), .O(n22999) );
  MAO222 U16992 ( .A1(n26344), .B1(gray_img[639]), .C1(n26343), .O(n26480) );
  MAO222S U16993 ( .A1(n26342), .B1(gray_img[638]), .C1(n26341), .O(n26343) );
  MAO222S U16994 ( .A1(n26340), .B1(gray_img[637]), .C1(n26339), .O(n26341) );
  MAO222 U16995 ( .A1(n26356), .B1(gray_img[631]), .C1(n26355), .O(n26360) );
  MAO222 U16996 ( .A1(n26354), .B1(gray_img[630]), .C1(n26353), .O(n26355) );
  MAO222 U16997 ( .A1(n26352), .B1(gray_img[629]), .C1(n26351), .O(n26353) );
  MAO222 U16998 ( .A1(n26204), .B1(n26203), .C1(n26202), .O(n26207) );
  MAO222S U16999 ( .A1(n26201), .B1(n26208), .C1(n26205), .O(n26204) );
  MAO222 U17000 ( .A1(n27053), .B1(n27051), .C1(n27043), .O(n27044) );
  MAO222 U17001 ( .A1(n27087), .B1(n27085), .C1(n27042), .O(n27043) );
  MAO222 U17002 ( .A1(n27092), .B1(n27090), .C1(n27041), .O(n27042) );
  MAO222 U17003 ( .A1(n27146), .B1(gray_img[583]), .C1(n27145), .O(n27159) );
  MAO222 U17004 ( .A1(n27144), .B1(gray_img[582]), .C1(n27143), .O(n27145) );
  MAO222 U17005 ( .A1(n27142), .B1(gray_img[581]), .C1(n27141), .O(n27143) );
  MAO222 U17006 ( .A1(n27140), .B1(gray_img[580]), .C1(n27139), .O(n27141) );
  MAO222 U17007 ( .A1(n27158), .B1(gray_img[591]), .C1(n27157), .O(n27244) );
  MAO222 U17008 ( .A1(n27156), .B1(gray_img[590]), .C1(n27155), .O(n27157) );
  MAO222 U17009 ( .A1(n27154), .B1(gray_img[589]), .C1(n27153), .O(n27155) );
  MAO222 U17010 ( .A1(n27167), .B1(n27166), .C1(n27165), .O(n27168) );
  MAO222S U17011 ( .A1(n27170), .B1(n27174), .C1(n27164), .O(n27165) );
  MAO222S U17012 ( .A1(n27202), .B1(n27206), .C1(n27163), .O(n27164) );
  MAO222S U17013 ( .A1(n27207), .B1(n27211), .C1(n27162), .O(n27163) );
  MAO222 U17014 ( .A1(n27622), .B1(gray_img[383]), .C1(n27621), .O(n27623) );
  MAO222S U17015 ( .A1(n27620), .B1(gray_img[382]), .C1(n27619), .O(n27621) );
  MAO222S U17016 ( .A1(n27618), .B1(gray_img[381]), .C1(n27617), .O(n27619) );
  MAO222S U17017 ( .A1(n27610), .B1(gray_img[375]), .C1(n27609), .O(n27657) );
  MAO222 U17018 ( .A1(n27608), .B1(gray_img[374]), .C1(n27607), .O(n27609) );
  MAO222S U17019 ( .A1(n27629), .B1(n27628), .C1(n15958), .O(n27631) );
  AO22S U17020 ( .A1(n27634), .A2(n27636), .B1(n27627), .B2(n15962), .O(n15958) );
  OR2S U17021 ( .I1(n27634), .I2(n27636), .O(n15962) );
  MAO222 U17022 ( .A1(n27641), .B1(n27639), .C1(n15957), .O(n27627) );
  MAO222 U17023 ( .A1(n27475), .B1(gray_img[359]), .C1(n27474), .O(n27776) );
  MAO222 U17024 ( .A1(n27473), .B1(gray_img[358]), .C1(n27472), .O(n27474) );
  MAO222 U17025 ( .A1(n27463), .B1(gray_img[495]), .C1(n27462), .O(n27476) );
  MAO222 U17026 ( .A1(n27461), .B1(gray_img[494]), .C1(n27460), .O(n27462) );
  MAO222S U17027 ( .A1(n27459), .B1(gray_img[493]), .C1(n27458), .O(n27460) );
  MAO222 U17028 ( .A1(n27484), .B1(n27483), .C1(n27482), .O(n27486) );
  MAO222S U17029 ( .A1(n27491), .B1(n27489), .C1(n27481), .O(n27482) );
  MAO222 U17030 ( .A1(n27496), .B1(n27494), .C1(n27480), .O(n27481) );
  MAO222 U17031 ( .A1(n27501), .B1(n27499), .C1(n27479), .O(n27480) );
  MAO222 U17032 ( .A1(gray_img[471]), .B1(n26774), .C1(n26773), .O(n26787) );
  MAO222S U17033 ( .A1(gray_img[470]), .B1(n26772), .C1(n26771), .O(n26773) );
  MAO222 U17034 ( .A1(n26784), .B1(gray_img[350]), .C1(n26783), .O(n26785) );
  MAO222S U17035 ( .A1(n26782), .B1(gray_img[349]), .C1(n26781), .O(n26783) );
  MAO222 U17036 ( .A1(n26795), .B1(n26794), .C1(n26793), .O(n26796) );
  MAO222 U17037 ( .A1(n26798), .B1(n26802), .C1(n26792), .O(n26793) );
  MAO222 U17038 ( .A1(n26803), .B1(n26807), .C1(n26791), .O(n26792) );
  MAO222S U17039 ( .A1(n26808), .B1(n26812), .C1(n26790), .O(n26791) );
  MAO222 U17040 ( .A1(n23387), .B1(gray_img[327]), .C1(n23386), .O(n23401) );
  MAO222 U17041 ( .A1(n23385), .B1(gray_img[326]), .C1(n23384), .O(n23386) );
  MAO222S U17042 ( .A1(n23400), .B1(gray_img[335]), .C1(n23399), .O(n23410) );
  MAO222 U17043 ( .A1(n23398), .B1(gray_img[334]), .C1(n23397), .O(n23399) );
  MAO222 U17044 ( .A1(n23396), .B1(gray_img[333]), .C1(n23395), .O(n23397) );
  MAO222S U17045 ( .A1(n27591), .B1(n27590), .C1(n27589), .O(n27593) );
  MAO222 U17046 ( .A1(n27420), .B1(gray_img[231]), .C1(n27419), .O(n27547) );
  MAO222 U17047 ( .A1(n27418), .B1(gray_img[230]), .C1(n27417), .O(n27419) );
  MOAI1S U17048 ( .A1(n27408), .A2(n27407), .B1(gray_img[111]), .B2(n27406), 
        .O(n27421) );
  MAO222S U17049 ( .A1(n27429), .B1(n27428), .C1(n27427), .O(n27431) );
  MAO222 U17050 ( .A1(n27436), .B1(n27434), .C1(n27426), .O(n27427) );
  MAO222 U17051 ( .A1(n27522), .B1(n27520), .C1(n27425), .O(n27426) );
  MAO222 U17052 ( .A1(n27527), .B1(n27525), .C1(n27424), .O(n27425) );
  MAO222 U17053 ( .A1(n16037), .B1(gray_img[87]), .C1(n16036), .O(n23483) );
  MAO222 U17054 ( .A1(n16035), .B1(gray_img[86]), .C1(n16034), .O(n16036) );
  MAO222S U17055 ( .A1(n16033), .B1(gray_img[85]), .C1(n16032), .O(n16034) );
  NR2 U17056 ( .I1(n16024), .I2(n16023), .O(n16038) );
  MAO222S U17057 ( .A1(gray_img[222]), .B1(n21141), .C1(n16021), .O(n16022) );
  MAO222S U17058 ( .A1(n20977), .B1(n20978), .C1(n15960), .O(n16044) );
  AO22S U17059 ( .A1(n26729), .A2(n26731), .B1(n16043), .B2(n15974), .O(n15960) );
  OR2S U17060 ( .I1(n26729), .I2(n26731), .O(n15974) );
  MAO222 U17061 ( .A1(n26833), .B1(n26831), .C1(n15959), .O(n16043) );
  MAO222 U17062 ( .A1(gray_img[207]), .B1(n23601), .C1(n23600), .O(n23615) );
  MAO222 U17063 ( .A1(gray_img[206]), .B1(n23599), .C1(n23598), .O(n23600) );
  MAO222 U17064 ( .A1(gray_img[205]), .B1(n23597), .C1(n23596), .O(n23598) );
  MAO222S U17065 ( .A1(gray_img[204]), .B1(n23595), .C1(n23594), .O(n23596) );
  MAO222S U17066 ( .A1(n23614), .B1(gray_img[71]), .C1(n23613), .O(n23624) );
  MAO222 U17067 ( .A1(n23612), .B1(gray_img[70]), .C1(n23611), .O(n23613) );
  MAO222 U17068 ( .A1(n23610), .B1(gray_img[69]), .C1(n23609), .O(n23611) );
  MAO222S U17069 ( .A1(n25261), .B1(n25262), .C1(n23621), .O(n23622) );
  MAO222S U17070 ( .A1(n23632), .B1(n23636), .C1(n23620), .O(n23621) );
  MAO222 U17071 ( .A1(n26888), .B1(n26886), .C1(n23619), .O(n23620) );
  MAO222 U17072 ( .A1(n26893), .B1(n26891), .C1(n23618), .O(n23619) );
  MAO222 U17073 ( .A1(n24975), .B1(gray_img[2015]), .C1(n23258), .O(n23276) );
  MAO222 U17074 ( .A1(n23257), .B1(gray_img[2014]), .C1(n23256), .O(n23258) );
  MAO222S U17075 ( .A1(n23255), .B1(gray_img[2013]), .C1(n23254), .O(n23256)
         );
  MAO222S U17076 ( .A1(n24981), .B1(n24982), .C1(n23282), .O(n23284) );
  MAO222 U17077 ( .A1(n25482), .B1(n25480), .C1(n23281), .O(n23282) );
  MAO222 U17078 ( .A1(n25587), .B1(n25585), .C1(n23280), .O(n23281) );
  MAO222S U17079 ( .A1(n25592), .B1(n25590), .C1(n23279), .O(n23280) );
  MAO222 U17080 ( .A1(n23430), .B1(gray_img[143]), .C1(n23429), .O(n30111) );
  MAO222 U17081 ( .A1(n23428), .B1(gray_img[142]), .C1(n23427), .O(n23429) );
  MAO222 U17082 ( .A1(n23426), .B1(gray_img[141]), .C1(n23425), .O(n23427) );
  MAO222 U17083 ( .A1(gray_img[135]), .B1(n25118), .C1(n23443), .O(n23444) );
  MAO222 U17084 ( .A1(gray_img[134]), .B1(n23442), .C1(n23441), .O(n23443) );
  MAO222 U17085 ( .A1(gray_img[133]), .B1(n23440), .C1(n23439), .O(n23441) );
  MAO222S U17086 ( .A1(n25113), .B1(n25114), .C1(n23449), .O(n23450) );
  MAO222S U17087 ( .A1(n23473), .B1(n23477), .C1(n23448), .O(n23449) );
  MAO222 U17088 ( .A1(n23468), .B1(n23472), .C1(n23447), .O(n23448) );
  MAO222 U17089 ( .A1(n23452), .B1(n23457), .C1(n15970), .O(n23447) );
  MUX2S U17090 ( .A(gray_img[649]), .B(gray_img[521]), .S(n29930), .O(n29970)
         );
  MUX2S U17091 ( .A(gray_img[929]), .B(gray_img[801]), .S(n28804), .O(n23241)
         );
  MUX2S U17092 ( .A(gray_img[457]), .B(gray_img[329]), .S(n23410), .O(n26938)
         );
  MUX2S U17093 ( .A(gray_img[592]), .B(gray_img[720]), .S(n27038), .O(n27113)
         );
  MUX2S U17094 ( .A(gray_img[593]), .B(gray_img[721]), .S(n27038), .O(n27120)
         );
  MUX2S U17095 ( .A(gray_img[233]), .B(gray_img[105]), .S(n27421), .O(n27542)
         );
  MUX2S U17096 ( .A(gray_img[648]), .B(gray_img[520]), .S(n29930), .O(n30011)
         );
  MUX2S U17097 ( .A(gray_img[1513]), .B(gray_img[1385]), .S(n28003), .O(n28133) );
  MUX2S U17098 ( .A(gray_img[1448]), .B(gray_img[1320]), .S(n28975), .O(n29016) );
  MUX2S U17099 ( .A(gray_img[1240]), .B(gray_img[1112]), .S(n28315), .O(n28431) );
  MUX2S U17100 ( .A(gray_img[1449]), .B(gray_img[1321]), .S(n28975), .O(n29039) );
  MUX2S U17101 ( .A(gray_img[905]), .B(gray_img[777]), .S(n29629), .O(n30017)
         );
  MUX2S U17102 ( .A(gray_img[880]), .B(gray_img[1008]), .S(n26401), .O(n26444)
         );
  MUX2S U17103 ( .A(gray_img[1241]), .B(gray_img[1113]), .S(n28315), .O(n28458) );
  MUX2S U17104 ( .A(gray_img[1881]), .B(gray_img[2009]), .S(n23276), .O(n25618) );
  MUX2S U17105 ( .A(gray_img[881]), .B(gray_img[1009]), .S(n26401), .O(n26472)
         );
  MUX2S U17106 ( .A(gray_img[545]), .B(gray_img[673]), .S(n28679), .O(n28705)
         );
  MUX2S U17107 ( .A(gray_img[753]), .B(gray_img[625]), .S(n26360), .O(n26478)
         );
  MUX2S U17108 ( .A(gray_img[1929]), .B(gray_img[1801]), .S(n29415), .O(n29492) );
  MUX2S U17109 ( .A(gray_img[161]), .B(gray_img[33]), .S(n26969), .O(n27377)
         );
  MUX2S U17110 ( .A(gray_img[1]), .B(gray_img[129]), .S(n23444), .O(n23478) );
  MUX2S U17111 ( .A(gray_img[1961]), .B(gray_img[1833]), .S(n30018), .O(n29193) );
  MUX2S U17112 ( .A(gray_img[1273]), .B(gray_img[1145]), .S(n23490), .O(n23367) );
  MUX2S U17113 ( .A(gray_img[857]), .B(gray_img[985]), .S(n23088), .O(n23120)
         );
  MAO222S U17114 ( .A1(n26183), .B1(gray_img[751]), .C1(n26182), .O(n26325) );
  MAO222 U17115 ( .A1(n26181), .B1(gray_img[750]), .C1(n26180), .O(n26182) );
  MAO222 U17116 ( .A1(n25537), .B1(gray_img[1759]), .C1(n25536), .O(n25577) );
  MAO222 U17117 ( .A1(n25535), .B1(gray_img[1758]), .C1(n25534), .O(n25536) );
  MAO222 U17118 ( .A1(n25533), .B1(gray_img[1757]), .C1(n25532), .O(n25534) );
  MAO222S U17119 ( .A1(n26639), .B1(gray_img[1031]), .C1(n26638), .O(n29731)
         );
  MAO222S U17120 ( .A1(n26637), .B1(gray_img[1030]), .C1(n26636), .O(n26638)
         );
  MAO222 U17121 ( .A1(n26635), .B1(gray_img[1029]), .C1(n26634), .O(n26636) );
  MUX2S U17122 ( .A(gray_img[1194]), .B(gray_img[1066]), .S(n29041), .O(n23044) );
  MUX2S U17123 ( .A(gray_img[1193]), .B(gray_img[1065]), .S(n29041), .O(n23372) );
  ND2S U17124 ( .I1(n25035), .I2(n25034), .O(n25047) );
  INV2 U17125 ( .I(cnt_cro_3b3[1]), .O(n24948) );
  OR2S U17126 ( .I1(n30360), .I2(n24945), .O(n24949) );
  ND2S U17127 ( .I1(n24945), .I2(n24948), .O(n24950) );
  OR2S U17128 ( .I1(n30438), .I2(n30440), .O(n15952) );
  MAO222S U17129 ( .A1(gray_scale_1[1]), .B1(n30435), .C1(gray_scale_1[0]), 
        .O(n19951) );
  ND3S U17130 ( .I1(n24955), .I2(n25040), .I3(cnt_cro_x[0]), .O(n24962) );
  ND2S U17131 ( .I1(cnt_bdyn[2]), .I2(n30302), .O(n30364) );
  ND2S U17132 ( .I1(n24942), .I2(n30359), .O(n30371) );
  ND3S U17133 ( .I1(n25041), .I2(n25040), .I3(cnt_cro_y[0]), .O(n25046) );
  NR2 U17134 ( .I1(n30411), .I2(n30255), .O(n24942) );
  INV1S U17135 ( .I(n24942), .O(n30360) );
  ND3S U17136 ( .I1(n21881), .I2(n21880), .I3(n21879), .O(n21882) );
  MAO222 U17137 ( .A1(n28746), .B1(gray_img[279]), .C1(n28745), .O(n28814) );
  MAO222 U17138 ( .A1(n28744), .B1(gray_img[278]), .C1(n28743), .O(n28745) );
  MAO222S U17139 ( .A1(n28742), .B1(gray_img[277]), .C1(n28741), .O(n28743) );
  MAO222S U17140 ( .A1(n28740), .B1(gray_img[276]), .C1(n28739), .O(n28741) );
  MAO222 U17141 ( .A1(n26123), .B1(gray_img[831]), .C1(n26122), .O(n28725) );
  MAO222 U17142 ( .A1(n26121), .B1(gray_img[830]), .C1(n26120), .O(n26122) );
  MAO222 U17143 ( .A1(n26119), .B1(gray_img[829]), .C1(n26118), .O(n26120) );
  MUX2S U17144 ( .A(gray_img[2016]), .B(gray_img[1888]), .S(n25861), .O(n26095) );
  MUX2S U17145 ( .A(gray_img[1880]), .B(gray_img[2008]), .S(n23276), .O(n23293) );
  MAO222 U17146 ( .A1(n26681), .B1(gray_img[1839]), .C1(n26680), .O(n30018) );
  MAO222 U17147 ( .A1(n26679), .B1(gray_img[1838]), .C1(n26678), .O(n26680) );
  MAO222 U17148 ( .A1(n26677), .B1(gray_img[1837]), .C1(n26676), .O(n26678) );
  MAO222 U17149 ( .A1(n26675), .B1(gray_img[1836]), .C1(n26674), .O(n26676) );
  MUX2S U17150 ( .A(gray_img[904]), .B(gray_img[776]), .S(n29629), .O(n30108)
         );
  MUX2S U17151 ( .A(gray_img[1928]), .B(gray_img[1800]), .S(n29415), .O(n30097) );
  MUX2S U17152 ( .A(gray_img[1784]), .B(gray_img[1656]), .S(n26009), .O(n26052) );
  MUX2S U17153 ( .A(gray_img[1640]), .B(gray_img[1768]), .S(n25805), .O(n25907) );
  MUX2S U17154 ( .A(gray_img[1608]), .B(gray_img[1736]), .S(n25679), .O(n25749) );
  MUX2S U17155 ( .A(gray_img[1712]), .B(gray_img[1584]), .S(n29222), .O(n29265) );
  MUX2S U17156 ( .A(gray_img[1704]), .B(gray_img[1576]), .S(n29121), .O(n29191) );
  MAO222 U17157 ( .A1(n26558), .B1(gray_img[1559]), .C1(n26557), .O(n29577) );
  MAO222 U17158 ( .A1(n26556), .B1(gray_img[1558]), .C1(n26555), .O(n26557) );
  MAO222S U17159 ( .A1(n26554), .B1(gray_img[1557]), .C1(n26553), .O(n26555)
         );
  MAO222 U17160 ( .A1(n28169), .B1(gray_img[567]), .C1(n28168), .O(n28215) );
  MAO222 U17161 ( .A1(n28167), .B1(gray_img[566]), .C1(n28166), .O(n28168) );
  MAO222 U17162 ( .A1(n28165), .B1(gray_img[565]), .C1(n28164), .O(n28166) );
  MAO222S U17163 ( .A1(n27917), .B1(gray_img[1527]), .C1(n27916), .O(n28134)
         );
  MAO222 U17164 ( .A1(n27915), .B1(gray_img[1526]), .C1(n27914), .O(n27916) );
  MAO222 U17165 ( .A1(n27913), .B1(gray_img[1525]), .C1(n27912), .O(n27914) );
  MAO222 U17166 ( .A1(n27911), .B1(gray_img[1524]), .C1(n27910), .O(n27912) );
  MUX2S U17167 ( .A(gray_img[1512]), .B(gray_img[1384]), .S(n28003), .O(n28213) );
  MAO222 U17168 ( .A1(n28632), .B1(gray_img[679]), .C1(n28631), .O(n28679) );
  MAO222 U17169 ( .A1(n28630), .B1(gray_img[678]), .C1(n28629), .O(n28631) );
  MAO222 U17170 ( .A1(n28628), .B1(gray_img[677]), .C1(n28627), .O(n28629) );
  MAO222 U17171 ( .A1(n28626), .B1(gray_img[676]), .C1(n28625), .O(n28627) );
  MUX2S U17172 ( .A(gray_img[1368]), .B(gray_img[1496]), .S(n28385), .O(n28606) );
  MAO222S U17173 ( .A1(n25199), .B1(gray_img[1359]), .C1(n23525), .O(n23536)
         );
  MAO222 U17174 ( .A1(n23524), .B1(gray_img[1358]), .C1(n23523), .O(n23525) );
  MAO222 U17175 ( .A1(n23522), .B1(gray_img[1357]), .C1(n23521), .O(n23523) );
  MUX2S U17176 ( .A(gray_img[528]), .B(gray_img[656]), .S(n29081), .O(n29358)
         );
  MUX2S U17177 ( .A(gray_img[1456]), .B(gray_img[1328]), .S(n18084), .O(n29349) );
  MUX2S U17178 ( .A(gray_img[1296]), .B(gray_img[1424]), .S(n29773), .O(n29903) );
  MAO222S U17179 ( .A1(n29668), .B1(gray_img[1423]), .C1(n29667), .O(n29991)
         );
  MAO222 U17180 ( .A1(n29666), .B1(gray_img[1422]), .C1(n29665), .O(n29667) );
  MAO222 U17181 ( .A1(n29664), .B1(gray_img[1421]), .C1(n29663), .O(n29665) );
  MAO222 U17182 ( .A1(n28506), .B1(gray_img[1095]), .C1(n28505), .O(n28669) );
  MAO222S U17183 ( .A1(n28504), .B1(gray_img[1094]), .C1(n28503), .O(n28505)
         );
  MAO222 U17184 ( .A1(n28502), .B1(gray_img[1093]), .C1(n28501), .O(n28503) );
  MUX2S U17185 ( .A(gray_img[1208]), .B(gray_img[1080]), .S(n28879), .O(n28942) );
  MUX2S U17186 ( .A(gray_img[152]), .B(gray_img[24]), .S(n27877), .O(n30086)
         );
  MUX2S U17187 ( .A(gray_img[312]), .B(gray_img[440]), .S(n26514), .O(n27850)
         );
  MUX2S U17188 ( .A(gray_img[1000]), .B(gray_img[872]), .S(n26256), .O(n27839)
         );
  MUX2S U17189 ( .A(gray_img[288]), .B(gray_img[416]), .S(n27288), .O(n30075)
         );
  MUX2S U17190 ( .A(n22990), .B(n30457), .S(n22994), .O(n23299) );
  MUX2S U17191 ( .A(gray_img[752]), .B(gray_img[624]), .S(n26360), .O(n26488)
         );
  MUX2S U17192 ( .A(gray_img[56]), .B(gray_img[184]), .S(n27735), .O(n27793)
         );
  MUX2S U17193 ( .A(gray_img[360]), .B(gray_img[488]), .S(n27476), .O(n27784)
         );
  MUX2S U17194 ( .A(gray_img[232]), .B(gray_img[104]), .S(n27421), .O(n27555)
         );
  OR2S U17195 ( .I1(n24652), .I2(n24693), .O(n24657) );
  OR2S U17196 ( .I1(n24653), .I2(n24695), .O(n24656) );
  ND3S U17197 ( .I1(n22045), .I2(n22044), .I3(n22043), .O(n22101) );
  ND3S U17198 ( .I1(n22155), .I2(n22154), .I3(n22153), .O(n22215) );
  MUX2S U17199 ( .A(gray_img[401]), .B(gray_img[273]), .S(n28814), .O(n28846)
         );
  MUX2S U17200 ( .A(gray_img[2033]), .B(gray_img[1905]), .S(n25970), .O(n26085) );
  MUX2S U17201 ( .A(gray_img[2017]), .B(gray_img[1889]), .S(n25861), .O(n25941) );
  MUX2S U17202 ( .A(gray_img[1993]), .B(gray_img[1865]), .S(n23582), .O(n25757) );
  MUX2S U17203 ( .A(gray_img[385]), .B(gray_img[257]), .S(n23360), .O(n30127)
         );
  MUX2S U17204 ( .A(gray_img[1785]), .B(gray_img[1657]), .S(n26009), .O(n26079) );
  MUX2S U17205 ( .A(gray_img[1609]), .B(gray_img[1737]), .S(n25679), .O(n25719) );
  MUX2S U17206 ( .A(gray_img[1713]), .B(gray_img[1585]), .S(n29222), .O(n29272) );
  MUX2S U17207 ( .A(gray_img[1705]), .B(gray_img[1577]), .S(n29121), .O(n29161) );
  MUX2S U17208 ( .A(gray_img[689]), .B(gray_img[561]), .S(n28215), .O(n28236)
         );
  MUX2S U17209 ( .A(gray_img[1393]), .B(gray_img[1521]), .S(n28134), .O(n27954) );
  MUX2S U17210 ( .A(gray_img[529]), .B(gray_img[657]), .S(n29081), .O(n29380)
         );
  MUX2S U17211 ( .A(gray_img[153]), .B(gray_img[25]), .S(n27877), .O(n28852)
         );
  MUX2S U17212 ( .A(gray_img[313]), .B(gray_img[441]), .S(n26514), .O(n27826)
         );
  MUX2S U17213 ( .A(gray_img[289]), .B(gray_img[417]), .S(n27288), .O(n27329)
         );
  MUX2S U17214 ( .A(gray_img[57]), .B(gray_img[185]), .S(n27735), .O(n27820)
         );
  MUX2S U17215 ( .A(gray_img[1297]), .B(gray_img[1425]), .S(n29773), .O(n29893) );
  MUX2S U17216 ( .A(gray_img[1169]), .B(gray_img[1041]), .S(n29853), .O(n29879) );
  MUX2S U17217 ( .A(gray_img[1001]), .B(gray_img[873]), .S(n26256), .O(n26296)
         );
  MUX2S U17218 ( .A(intadd_99_CI), .B(n22989), .S(n22994), .O(n27229) );
  MUX2S U17219 ( .A(gray_img[969]), .B(gray_img[841]), .S(n23295), .O(n27225)
         );
  MUX2S U17220 ( .A(gray_img[713]), .B(gray_img[585]), .S(n27244), .O(n27250)
         );
  MUX2S U17221 ( .A(gray_img[361]), .B(gray_img[489]), .S(n27476), .O(n27517)
         );
  AOI12HS U17222 ( .B1(mem_data_a_out[1]), .B2(n16010), .A1(n18475), .O(n29884) );
  MUX2S U17223 ( .A(gray_img[193]), .B(gray_img[65]), .S(n23624), .O(n26930)
         );
  MUX2S U17224 ( .A(gray_img[1457]), .B(gray_img[1329]), .S(n18084), .O(n28919) );
  ND3S U17225 ( .I1(n22484), .I2(n22483), .I3(n22482), .O(n22539) );
  ND3S U17226 ( .I1(n22594), .I2(n22593), .I3(n22592), .O(n22653) );
  MUX2S U17227 ( .A(gray_img[402]), .B(gray_img[274]), .S(n28814), .O(n28800)
         );
  MUX2S U17228 ( .A(gray_img[954]), .B(gray_img[826]), .S(n28725), .O(n28231)
         );
  MUX2S U17229 ( .A(gray_img[2034]), .B(gray_img[1906]), .S(n25970), .O(n26072) );
  MUX2S U17230 ( .A(gray_img[2018]), .B(gray_img[1890]), .S(n25861), .O(n25927) );
  MUX2S U17231 ( .A(gray_img[930]), .B(gray_img[802]), .S(n28804), .O(n28700)
         );
  MUX2S U17232 ( .A(gray_img[1882]), .B(gray_img[2010]), .S(n23276), .O(n25602) );
  MUX2S U17233 ( .A(gray_img[1994]), .B(gray_img[1866]), .S(n23582), .O(n25739) );
  MUX2S U17234 ( .A(gray_img[386]), .B(gray_img[258]), .S(n23360), .O(n30062)
         );
  MUX2S U17235 ( .A(gray_img[922]), .B(gray_img[794]), .S(n29299), .O(n29373)
         );
  MUX2S U17236 ( .A(gray_img[1962]), .B(gray_img[1834]), .S(n30018), .O(n29177) );
  MUX2S U17237 ( .A(gray_img[906]), .B(gray_img[778]), .S(n29629), .O(n29990)
         );
  MUX2S U17238 ( .A(gray_img[1946]), .B(gray_img[1818]), .S(n29517), .O(n29576) );
  MUX2S U17239 ( .A(gray_img[1930]), .B(gray_img[1802]), .S(n29415), .O(n29476) );
  MUX2S U17240 ( .A(gray_img[1786]), .B(gray_img[1658]), .S(n26009), .O(n26044) );
  MUX2S U17241 ( .A(gray_img[1642]), .B(gray_img[1770]), .S(n25805), .O(n25896) );
  MUX2S U17242 ( .A(gray_img[1610]), .B(gray_img[1738]), .S(n25679), .O(n25714) );
  MUX2S U17243 ( .A(gray_img[1714]), .B(gray_img[1586]), .S(n29222), .O(n29257) );
  MUX2S U17244 ( .A(gray_img[1706]), .B(gray_img[1578]), .S(n29121), .O(n29156) );
  MUX2S U17245 ( .A(gray_img[690]), .B(gray_img[562]), .S(n28215), .O(n28196)
         );
  MUX2S U17246 ( .A(gray_img[1394]), .B(gray_img[1522]), .S(n28134), .O(n27949) );
  MUX2S U17247 ( .A(gray_img[1514]), .B(gray_img[1386]), .S(n28003), .O(n28120) );
  MUX2S U17248 ( .A(gray_img[546]), .B(gray_img[674]), .S(n28679), .O(n28664)
         );
  MUX2S U17249 ( .A(gray_img[530]), .B(gray_img[658]), .S(n29081), .O(n29339)
         );
  MUX2S U17250 ( .A(gray_img[650]), .B(gray_img[522]), .S(n29930), .O(n29965)
         );
  MUX2S U17251 ( .A(gray_img[154]), .B(gray_img[26]), .S(n27877), .O(n28839)
         );
  MUX2S U17252 ( .A(gray_img[314]), .B(gray_img[442]), .S(n26514), .O(n27813)
         );
  MUX2S U17253 ( .A(gray_img[290]), .B(gray_img[418]), .S(n27288), .O(n27324)
         );
  MUX2S U17254 ( .A(gray_img[58]), .B(gray_img[186]), .S(n27735), .O(n27771)
         );
  MUX2S U17255 ( .A(gray_img[162]), .B(gray_img[34]), .S(n26969), .O(n27349)
         );
  MUX2S U17256 ( .A(gray_img[1458]), .B(gray_img[1330]), .S(n18084), .O(n28914) );
  MUX2S U17257 ( .A(gray_img[1450]), .B(gray_img[1322]), .S(n28975), .O(n29008) );
  MUX2S U17258 ( .A(gray_img[1298]), .B(gray_img[1426]), .S(n29773), .O(n29878) );
  MUX2S U17259 ( .A(gray_img[1290]), .B(gray_img[1418]), .S(n29991), .O(n29701) );
  MUX2S U17260 ( .A(gray_img[1274]), .B(gray_img[1146]), .S(n23490), .O(n23335) );
  MUX2S U17261 ( .A(gray_img[1242]), .B(gray_img[1114]), .S(n28315), .O(n28420) );
  MUX2S U17262 ( .A(gray_img[1218]), .B(gray_img[1090]), .S(n28669), .O(n28576) );
  MUX2S U17263 ( .A(gray_img[1210]), .B(gray_img[1082]), .S(n28879), .O(n28934) );
  MUX2S U17264 ( .A(gray_img[1170]), .B(gray_img[1042]), .S(n29853), .O(n29847) );
  MUX2S U17265 ( .A(gray_img[1154]), .B(gray_img[1026]), .S(n29731), .O(n29726) );
  MUX2S U17266 ( .A(gray_img[882]), .B(gray_img[1010]), .S(n26401), .O(n26436)
         );
  MUX2S U17267 ( .A(gray_img[1002]), .B(gray_img[874]), .S(n26256), .O(n26291)
         );
  MUX2S U17268 ( .A(gray_img[858]), .B(gray_img[986]), .S(n23088), .O(n23095)
         );
  MUX2S U17269 ( .A(n22988), .B(n22987), .S(n22994), .O(n27221) );
  MUX2S U17270 ( .A(gray_img[970]), .B(gray_img[842]), .S(n23295), .O(n27218)
         );
  MUX2S U17271 ( .A(gray_img[754]), .B(gray_img[626]), .S(n26360), .O(n26465)
         );
  MUX2S U17272 ( .A(gray_img[594]), .B(gray_img[722]), .S(n27038), .O(n27102)
         );
  MUX2S U17273 ( .A(gray_img[714]), .B(gray_img[586]), .S(n27244), .O(n27236)
         );
  MUX2S U17274 ( .A(gray_img[506]), .B(gray_img[378]), .S(n27623), .O(n27656)
         );
  MUX2S U17275 ( .A(gray_img[362]), .B(gray_img[490]), .S(n27476), .O(n27511)
         );
  MUX2S U17276 ( .A(gray_img[474]), .B(gray_img[346]), .S(n27353), .O(n26818)
         );
  MUX2S U17277 ( .A(gray_img[458]), .B(gray_img[330]), .S(n23410), .O(n26923)
         );
  MUX2S U17278 ( .A(gray_img[242]), .B(gray_img[114]), .S(n27586), .O(n27684)
         );
  MUX2S U17279 ( .A(gray_img[234]), .B(gray_img[106]), .S(n27421), .O(n27537)
         );
  MUX2S U17280 ( .A(gray_img[194]), .B(gray_img[66]), .S(n23624), .O(n26903)
         );
  MUX2S U17281 ( .A(gray_img[1370]), .B(gray_img[1498]), .S(n28385), .O(n28451) );
  ND3S U17282 ( .I1(n22324), .I2(n22323), .I3(n22322), .O(n22325) );
  ND3S U17283 ( .I1(n22272), .I2(n22271), .I3(n22270), .O(n22326) );
  MUX2S U17284 ( .A(gray_img[2]), .B(gray_img[130]), .S(n23444), .O(n23463) );
  AOI12HS U17285 ( .B1(mem_data_a_out[2]), .B2(n16010), .A1(n18483), .O(n29849) );
  MUX2S U17286 ( .A(gray_img[403]), .B(gray_img[275]), .S(n28814), .O(n28795)
         );
  MUX2S U17287 ( .A(gray_img[955]), .B(gray_img[827]), .S(n28725), .O(n28226)
         );
  MUX2S U17288 ( .A(gray_img[2035]), .B(gray_img[1907]), .S(n25970), .O(n26067) );
  MUX2S U17289 ( .A(gray_img[2019]), .B(gray_img[1891]), .S(n25861), .O(n25922) );
  MUX2S U17290 ( .A(gray_img[931]), .B(gray_img[803]), .S(n28804), .O(n28695)
         );
  MUX2S U17291 ( .A(gray_img[1883]), .B(gray_img[2011]), .S(n23276), .O(n25597) );
  MUX2S U17292 ( .A(gray_img[1995]), .B(gray_img[1867]), .S(n23582), .O(n25734) );
  MUX2S U17293 ( .A(gray_img[387]), .B(gray_img[259]), .S(n23360), .O(n30055)
         );
  MUX2S U17294 ( .A(gray_img[923]), .B(gray_img[795]), .S(n29299), .O(n29368)
         );
  MUX2S U17295 ( .A(gray_img[1971]), .B(gray_img[1843]), .S(n23162), .O(n23168) );
  MUX2S U17296 ( .A(gray_img[1963]), .B(gray_img[1835]), .S(n30018), .O(n29172) );
  MUX2S U17297 ( .A(gray_img[907]), .B(gray_img[779]), .S(n29629), .O(n29985)
         );
  MUX2S U17298 ( .A(gray_img[1947]), .B(gray_img[1819]), .S(n29517), .O(n29571) );
  MUX2S U17299 ( .A(gray_img[1931]), .B(gray_img[1803]), .S(n29415), .O(n29471) );
  MUX2S U17300 ( .A(gray_img[1787]), .B(gray_img[1659]), .S(n26009), .O(n26039) );
  MUX2S U17301 ( .A(gray_img[1643]), .B(gray_img[1771]), .S(n25805), .O(n25891) );
  MUX2S U17302 ( .A(gray_img[1627]), .B(gray_img[1755]), .S(n25577), .O(n25564) );
  MUX2S U17303 ( .A(gray_img[1611]), .B(gray_img[1739]), .S(n25679), .O(n25709) );
  MUX2S U17304 ( .A(gray_img[1715]), .B(gray_img[1587]), .S(n29222), .O(n29252) );
  MUX2S U17305 ( .A(gray_img[1707]), .B(gray_img[1579]), .S(n29121), .O(n29151) );
  MUX2S U17306 ( .A(gray_img[1675]), .B(gray_img[1547]), .S(n26601), .O(n29446) );
  MUX2S U17307 ( .A(gray_img[691]), .B(gray_img[563]), .S(n28215), .O(n28191)
         );
  MUX2S U17308 ( .A(gray_img[547]), .B(gray_img[675]), .S(n28679), .O(n28659)
         );
  MUX2S U17309 ( .A(gray_img[531]), .B(gray_img[659]), .S(n29081), .O(n29334)
         );
  MUX2S U17310 ( .A(gray_img[651]), .B(gray_img[523]), .S(n29930), .O(n29960)
         );
  MUX2S U17311 ( .A(gray_img[155]), .B(gray_img[27]), .S(n27877), .O(n28834)
         );
  MUX2S U17312 ( .A(gray_img[315]), .B(gray_img[443]), .S(n26514), .O(n27808)
         );
  MUX2S U17313 ( .A(gray_img[291]), .B(gray_img[419]), .S(n27288), .O(n27319)
         );
  MUX2S U17314 ( .A(gray_img[59]), .B(gray_img[187]), .S(n27735), .O(n27766)
         );
  MUX2S U17315 ( .A(gray_img[163]), .B(gray_img[35]), .S(n26969), .O(n27344)
         );
  MUX2S U17316 ( .A(gray_img[1515]), .B(gray_img[1387]), .S(n28003), .O(n28115) );
  MUX2S U17317 ( .A(gray_img[1371]), .B(gray_img[1499]), .S(n28385), .O(n28446) );
  MUX2S U17318 ( .A(gray_img[1459]), .B(gray_img[1331]), .S(n18084), .O(n28909) );
  MUX2S U17319 ( .A(gray_img[1451]), .B(gray_img[1323]), .S(n28975), .O(n29003) );
  MUX2S U17320 ( .A(gray_img[1299]), .B(gray_img[1427]), .S(n29773), .O(n29873) );
  MUX2S U17321 ( .A(gray_img[1291]), .B(gray_img[1419]), .S(n29991), .O(n29696) );
  MUX2S U17322 ( .A(gray_img[1275]), .B(gray_img[1147]), .S(n23490), .O(n23345) );
  MUX2S U17323 ( .A(gray_img[1131]), .B(gray_img[1259]), .S(n28056), .O(n28084) );
  MUX2S U17324 ( .A(gray_img[1243]), .B(gray_img[1115]), .S(n28315), .O(n28415) );
  MUX2S U17325 ( .A(gray_img[1219]), .B(gray_img[1091]), .S(n28669), .O(n28571) );
  MUX2S U17326 ( .A(gray_img[1211]), .B(gray_img[1083]), .S(n28879), .O(n28929) );
  MUX2S U17327 ( .A(gray_img[1195]), .B(gray_img[1067]), .S(n29041), .O(n29027) );
  MUX2S U17328 ( .A(gray_img[1171]), .B(gray_img[1043]), .S(n29853), .O(n29841) );
  MUX2S U17329 ( .A(gray_img[1155]), .B(gray_img[1027]), .S(n29731), .O(n29721) );
  MUX2S U17330 ( .A(gray_img[883]), .B(gray_img[1011]), .S(n26401), .O(n26431)
         );
  MUX2S U17331 ( .A(gray_img[1003]), .B(gray_img[875]), .S(n26256), .O(n26286)
         );
  MUX2S U17332 ( .A(gray_img[859]), .B(gray_img[987]), .S(n23088), .O(n23100)
         );
  MUX2S U17333 ( .A(n22986), .B(n22985), .S(n22994), .O(n27216) );
  MUX2S U17334 ( .A(gray_img[971]), .B(gray_img[843]), .S(n23295), .O(n27213)
         );
  MUX2S U17335 ( .A(gray_img[755]), .B(gray_img[627]), .S(n26360), .O(n26460)
         );
  MUX2S U17336 ( .A(gray_img[595]), .B(gray_img[723]), .S(n27038), .O(n27097)
         );
  MUX2S U17337 ( .A(gray_img[715]), .B(gray_img[587]), .S(n27244), .O(n27231)
         );
  MUX2S U17338 ( .A(gray_img[507]), .B(gray_img[379]), .S(n27623), .O(n27651)
         );
  MUX2S U17339 ( .A(gray_img[363]), .B(gray_img[491]), .S(n27476), .O(n27506)
         );
  MUX2S U17340 ( .A(gray_img[475]), .B(gray_img[347]), .S(n27353), .O(n26813)
         );
  MUX2S U17341 ( .A(gray_img[459]), .B(gray_img[331]), .S(n23410), .O(n26918)
         );
  MUX2S U17342 ( .A(gray_img[243]), .B(gray_img[115]), .S(n27586), .O(n27679)
         );
  MUX2S U17343 ( .A(gray_img[235]), .B(gray_img[107]), .S(n27421), .O(n27532)
         );
  MUX2S U17344 ( .A(gray_img[211]), .B(gray_img[83]), .S(n23483), .O(n16063)
         );
  MUX2S U17345 ( .A(gray_img[195]), .B(gray_img[67]), .S(n23624), .O(n26898)
         );
  MUX2S U17346 ( .A(gray_img[1395]), .B(gray_img[1523]), .S(n28134), .O(n27944) );
  ND3S U17347 ( .I1(n21449), .I2(n21448), .I3(n21447), .O(n21450) );
  ND3S U17348 ( .I1(n21399), .I2(n21398), .I3(n21397), .O(n21451) );
  MUX2S U17349 ( .A(gray_img[3]), .B(gray_img[131]), .S(n23444), .O(n23458) );
  AOI12HS U17350 ( .B1(mem_data_a_out[3]), .B2(n16010), .A1(n16065), .O(n29843) );
  MUX2S U17351 ( .A(gray_img[404]), .B(gray_img[276]), .S(n28814), .O(n28790)
         );
  MUX2S U17352 ( .A(gray_img[956]), .B(gray_img[828]), .S(n28725), .O(n28221)
         );
  MUX2S U17353 ( .A(gray_img[2036]), .B(gray_img[1908]), .S(n25970), .O(n26062) );
  MUX2S U17354 ( .A(gray_img[2020]), .B(gray_img[1892]), .S(n25861), .O(n25917) );
  MUX2S U17355 ( .A(gray_img[932]), .B(gray_img[804]), .S(n28804), .O(n28690)
         );
  MUX2S U17356 ( .A(gray_img[1884]), .B(gray_img[2012]), .S(n23276), .O(n25592) );
  MUX2S U17357 ( .A(gray_img[1996]), .B(gray_img[1868]), .S(n23582), .O(n25729) );
  MUX2S U17358 ( .A(gray_img[388]), .B(gray_img[260]), .S(n23360), .O(n30049)
         );
  MUX2S U17359 ( .A(gray_img[924]), .B(gray_img[796]), .S(n29299), .O(n29363)
         );
  MUX2S U17360 ( .A(gray_img[1964]), .B(gray_img[1836]), .S(n30018), .O(n29167) );
  MUX2S U17361 ( .A(gray_img[908]), .B(gray_img[780]), .S(n29629), .O(n29980)
         );
  MUX2S U17362 ( .A(gray_img[692]), .B(gray_img[564]), .S(n28215), .O(n28186)
         );
  MUX2S U17363 ( .A(gray_img[548]), .B(gray_img[676]), .S(n28679), .O(n28654)
         );
  MUX2S U17364 ( .A(gray_img[532]), .B(gray_img[660]), .S(n29081), .O(n29329)
         );
  MUX2S U17365 ( .A(gray_img[652]), .B(gray_img[524]), .S(n29930), .O(n29955)
         );
  MUX2S U17366 ( .A(gray_img[156]), .B(gray_img[28]), .S(n27877), .O(n28829)
         );
  MUX2S U17367 ( .A(gray_img[316]), .B(gray_img[444]), .S(n26514), .O(n27803)
         );
  MUX2S U17368 ( .A(gray_img[292]), .B(gray_img[420]), .S(n27288), .O(n27313)
         );
  MUX2S U17369 ( .A(gray_img[60]), .B(gray_img[188]), .S(n27735), .O(n27761)
         );
  MUX2S U17370 ( .A(gray_img[164]), .B(gray_img[36]), .S(n26969), .O(n27339)
         );
  MUX2S U17371 ( .A(gray_img[1932]), .B(gray_img[1804]), .S(n29415), .O(n29466) );
  MUX2S U17372 ( .A(gray_img[1788]), .B(gray_img[1660]), .S(n26009), .O(n26034) );
  MUX2S U17373 ( .A(gray_img[1644]), .B(gray_img[1772]), .S(n25805), .O(n25886) );
  MUX2S U17374 ( .A(gray_img[1612]), .B(gray_img[1740]), .S(n25679), .O(n25704) );
  MUX2S U17375 ( .A(gray_img[1716]), .B(gray_img[1588]), .S(n29222), .O(n29247) );
  MUX2S U17376 ( .A(gray_img[1708]), .B(gray_img[1580]), .S(n29121), .O(n29146) );
  MUX2S U17377 ( .A(gray_img[1676]), .B(gray_img[1548]), .S(n26601), .O(n29441) );
  MUX2S U17378 ( .A(gray_img[1396]), .B(gray_img[1524]), .S(n28134), .O(n27939) );
  MUX2S U17379 ( .A(gray_img[1516]), .B(gray_img[1388]), .S(n28003), .O(n28110) );
  MUX2S U17380 ( .A(gray_img[1372]), .B(gray_img[1500]), .S(n28385), .O(n28441) );
  MUX2S U17381 ( .A(gray_img[1460]), .B(gray_img[1332]), .S(n18084), .O(n23202) );
  MUX2S U17382 ( .A(gray_img[1452]), .B(gray_img[1324]), .S(n28975), .O(n28998) );
  MUX2S U17383 ( .A(gray_img[1300]), .B(gray_img[1428]), .S(n29773), .O(n29868) );
  MUX2S U17384 ( .A(gray_img[1292]), .B(gray_img[1420]), .S(n29991), .O(n29691) );
  MUX2S U17385 ( .A(gray_img[1276]), .B(gray_img[1148]), .S(n23490), .O(n23355) );
  MUX2S U17386 ( .A(gray_img[1132]), .B(gray_img[1260]), .S(n28056), .O(n28079) );
  MUX2S U17387 ( .A(gray_img[1244]), .B(gray_img[1116]), .S(n28315), .O(n28410) );
  MUX2S U17388 ( .A(gray_img[1220]), .B(gray_img[1092]), .S(n28669), .O(n28566) );
  MUX2S U17389 ( .A(gray_img[1212]), .B(gray_img[1084]), .S(n28879), .O(n28924) );
  MUX2S U17390 ( .A(gray_img[1196]), .B(gray_img[1068]), .S(n29041), .O(n29022) );
  MUX2S U17391 ( .A(gray_img[1172]), .B(gray_img[1044]), .S(n29853), .O(n29835) );
  MUX2S U17392 ( .A(gray_img[884]), .B(gray_img[1012]), .S(n26401), .O(n26426)
         );
  MUX2S U17393 ( .A(gray_img[1004]), .B(gray_img[876]), .S(n26256), .O(n26281)
         );
  MUX2S U17394 ( .A(gray_img[860]), .B(gray_img[988]), .S(n23088), .O(n23105)
         );
  MUX2S U17395 ( .A(n22984), .B(n22983), .S(n22994), .O(n27201) );
  MUX2S U17396 ( .A(gray_img[972]), .B(gray_img[844]), .S(n23295), .O(n27198)
         );
  MUX2S U17397 ( .A(gray_img[756]), .B(gray_img[628]), .S(n26360), .O(n26455)
         );
  MUX2S U17398 ( .A(gray_img[596]), .B(gray_img[724]), .S(n27038), .O(n27092)
         );
  MUX2S U17399 ( .A(gray_img[716]), .B(gray_img[588]), .S(n27244), .O(n27207)
         );
  MUX2S U17400 ( .A(gray_img[508]), .B(gray_img[380]), .S(n27623), .O(n27646)
         );
  MUX2S U17401 ( .A(gray_img[364]), .B(gray_img[492]), .S(n27476), .O(n27501)
         );
  MUX2S U17402 ( .A(gray_img[476]), .B(gray_img[348]), .S(n27353), .O(n26808)
         );
  MUX2S U17403 ( .A(gray_img[460]), .B(gray_img[332]), .S(n23410), .O(n26913)
         );
  MUX2S U17404 ( .A(gray_img[244]), .B(gray_img[116]), .S(n27586), .O(n27674)
         );
  MUX2S U17405 ( .A(gray_img[236]), .B(gray_img[108]), .S(n27421), .O(n27527)
         );
  MUX2S U17406 ( .A(gray_img[196]), .B(gray_img[68]), .S(n23624), .O(n26893)
         );
  MUX2S U17407 ( .A(gray_img[1948]), .B(gray_img[1820]), .S(n29517), .O(n29565) );
  ND3S U17408 ( .I1(n21721), .I2(n21720), .I3(n21719), .O(n21773) );
  ND3S U17409 ( .I1(n21662), .I2(n21661), .I3(n21660), .O(n21663) );
  MUX2S U17410 ( .A(gray_img[4]), .B(gray_img[132]), .S(n23444), .O(n23452) );
  MUX2S U17411 ( .A(gray_img[405]), .B(gray_img[277]), .S(n28814), .O(n28785)
         );
  MUX2S U17412 ( .A(gray_img[957]), .B(gray_img[829]), .S(n28725), .O(n28255)
         );
  MUX2S U17413 ( .A(gray_img[2037]), .B(gray_img[1909]), .S(n25970), .O(n26057) );
  MUX2S U17414 ( .A(gray_img[2021]), .B(gray_img[1893]), .S(n25861), .O(n25912) );
  MUX2S U17415 ( .A(gray_img[933]), .B(gray_img[805]), .S(n28804), .O(n28685)
         );
  MUX2S U17416 ( .A(gray_img[1885]), .B(gray_img[2013]), .S(n23276), .O(n25587) );
  MUX2S U17417 ( .A(gray_img[1997]), .B(gray_img[1869]), .S(n23582), .O(n25724) );
  MUX2S U17418 ( .A(gray_img[389]), .B(gray_img[261]), .S(n23360), .O(n30043)
         );
  MUX2S U17419 ( .A(gray_img[909]), .B(gray_img[781]), .S(n29629), .O(n29975)
         );
  MUX2S U17420 ( .A(gray_img[693]), .B(gray_img[565]), .S(n28215), .O(n28246)
         );
  MUX2S U17421 ( .A(gray_img[549]), .B(gray_img[677]), .S(n28679), .O(n28649)
         );
  MUX2S U17422 ( .A(gray_img[533]), .B(gray_img[661]), .S(n29081), .O(n29319)
         );
  MUX2S U17423 ( .A(gray_img[653]), .B(gray_img[525]), .S(n29930), .O(n29950)
         );
  MUX2S U17424 ( .A(gray_img[157]), .B(gray_img[29]), .S(n27877), .O(n28824)
         );
  MUX2S U17425 ( .A(gray_img[317]), .B(gray_img[445]), .S(n26514), .O(n27798)
         );
  MUX2S U17426 ( .A(gray_img[293]), .B(gray_img[421]), .S(n27288), .O(n27308)
         );
  MUX2S U17427 ( .A(gray_img[61]), .B(gray_img[189]), .S(n27735), .O(n27756)
         );
  MUX2S U17428 ( .A(gray_img[165]), .B(gray_img[37]), .S(n26969), .O(n27334)
         );
  MUX2S U17429 ( .A(gray_img[925]), .B(gray_img[797]), .S(n29299), .O(n29324)
         );
  MUX2S U17430 ( .A(gray_img[1965]), .B(gray_img[1837]), .S(n30018), .O(n29162) );
  MUX2S U17431 ( .A(gray_img[1949]), .B(gray_img[1821]), .S(n29517), .O(n29560) );
  MUX2S U17432 ( .A(gray_img[1933]), .B(gray_img[1805]), .S(n29415), .O(n29461) );
  MUX2S U17433 ( .A(gray_img[1789]), .B(gray_img[1661]), .S(n26009), .O(n26029) );
  MUX2S U17434 ( .A(gray_img[1645]), .B(gray_img[1773]), .S(n25805), .O(n25881) );
  MUX2S U17435 ( .A(gray_img[1629]), .B(gray_img[1757]), .S(n25577), .O(n25554) );
  MUX2S U17436 ( .A(gray_img[1613]), .B(gray_img[1741]), .S(n25679), .O(n25699) );
  MUX2S U17437 ( .A(gray_img[1717]), .B(gray_img[1589]), .S(n29222), .O(n29242) );
  MUX2S U17438 ( .A(gray_img[1709]), .B(gray_img[1581]), .S(n29121), .O(n29141) );
  MUX2S U17439 ( .A(gray_img[1677]), .B(gray_img[1549]), .S(n26601), .O(n29436) );
  MUX2S U17440 ( .A(gray_img[1397]), .B(gray_img[1525]), .S(n28134), .O(n27934) );
  MUX2S U17441 ( .A(gray_img[1517]), .B(gray_img[1389]), .S(n28003), .O(n28105) );
  MUX2S U17442 ( .A(gray_img[1373]), .B(gray_img[1501]), .S(n28385), .O(n28436) );
  MUX2S U17443 ( .A(gray_img[1485]), .B(gray_img[1357]), .S(n23536), .O(n28542) );
  MUX2S U17444 ( .A(gray_img[1461]), .B(gray_img[1333]), .S(n18084), .O(n28899) );
  MUX2S U17445 ( .A(gray_img[1453]), .B(gray_img[1325]), .S(n28975), .O(n28993) );
  MUX2S U17446 ( .A(gray_img[1301]), .B(gray_img[1429]), .S(n29773), .O(n29863) );
  MUX2S U17447 ( .A(gray_img[1293]), .B(gray_img[1421]), .S(n29991), .O(n29686) );
  MUX2S U17448 ( .A(gray_img[1277]), .B(gray_img[1149]), .S(n23490), .O(n23340) );
  MUX2S U17449 ( .A(gray_img[1133]), .B(gray_img[1261]), .S(n28056), .O(n28074) );
  MUX2S U17450 ( .A(gray_img[1245]), .B(gray_img[1117]), .S(n28315), .O(n28405) );
  MUX2S U17451 ( .A(gray_img[1221]), .B(gray_img[1093]), .S(n28669), .O(n28561) );
  MUX2S U17452 ( .A(gray_img[1213]), .B(gray_img[1085]), .S(n28879), .O(n28904) );
  MUX2S U17453 ( .A(gray_img[1197]), .B(gray_img[1069]), .S(n29041), .O(n29017) );
  MUX2S U17454 ( .A(gray_img[1173]), .B(gray_img[1045]), .S(n29853), .O(n29829) );
  MUX2S U17455 ( .A(gray_img[1157]), .B(gray_img[1029]), .S(n29731), .O(n29711) );
  MUX2S U17456 ( .A(gray_img[885]), .B(gray_img[1013]), .S(n26401), .O(n26421)
         );
  MUX2S U17457 ( .A(gray_img[1005]), .B(gray_img[877]), .S(n26256), .O(n26276)
         );
  MUX2S U17458 ( .A(gray_img[861]), .B(gray_img[989]), .S(n23088), .O(n23110)
         );
  MUX2S U17459 ( .A(gray_img[757]), .B(gray_img[629]), .S(n26360), .O(n26450)
         );
  ND2S U17460 ( .I1(n20930), .I2(n25374), .O(n26322) );
  MUX2S U17461 ( .A(gray_img[597]), .B(gray_img[725]), .S(n27038), .O(n27087)
         );
  MUX2S U17462 ( .A(gray_img[717]), .B(gray_img[589]), .S(n27244), .O(n27202)
         );
  MUX2S U17463 ( .A(gray_img[509]), .B(gray_img[381]), .S(n27623), .O(n27641)
         );
  MUX2S U17464 ( .A(gray_img[365]), .B(gray_img[493]), .S(n27476), .O(n27496)
         );
  MUX2S U17465 ( .A(gray_img[461]), .B(gray_img[333]), .S(n23410), .O(n26908)
         );
  MUX2S U17466 ( .A(gray_img[245]), .B(gray_img[117]), .S(n27586), .O(n27669)
         );
  MUX2S U17467 ( .A(gray_img[237]), .B(gray_img[109]), .S(n27421), .O(n27522)
         );
  MUX2S U17468 ( .A(gray_img[213]), .B(gray_img[85]), .S(n23483), .O(n26833)
         );
  MUX2S U17469 ( .A(gray_img[197]), .B(gray_img[69]), .S(n23624), .O(n26888)
         );
  ND3S U17470 ( .I1(n22955), .I2(n22954), .I3(n22953), .O(n22956) );
  ND3S U17471 ( .I1(n22717), .I2(n22716), .I3(n22715), .O(n22783) );
  MUX2S U17472 ( .A(gray_img[5]), .B(gray_img[133]), .S(n23444), .O(n23468) );
  MUX2S U17473 ( .A(gray_img[406]), .B(gray_img[278]), .S(n28814), .O(n28780)
         );
  ND2S U17474 ( .I1(n20918), .I2(n25374), .O(n28840) );
  NR2 U17475 ( .I1(n29680), .I2(n26134), .O(n28727) );
  INV1S U17476 ( .I(n26133), .O(n26134) );
  MUX2S U17477 ( .A(gray_img[958]), .B(gray_img[830]), .S(n28725), .O(n26135)
         );
  ND2S U17478 ( .I1(n20884), .I2(n25374), .O(n28728) );
  OR2 U17479 ( .I1(n29680), .I2(n26133), .O(n28733) );
  MUX2S U17480 ( .A(gray_img[2038]), .B(gray_img[1910]), .S(n25970), .O(n25983) );
  ND2S U17481 ( .I1(n21065), .I2(n25374), .O(n28718) );
  MUX2S U17482 ( .A(gray_img[2022]), .B(gray_img[1894]), .S(n25861), .O(n25876) );
  ND2S U17483 ( .I1(n25075), .I2(n25374), .O(n26090) );
  ND2S U17484 ( .I1(n23242), .I2(n25374), .O(n28807) );
  INV1S U17485 ( .I(n23239), .O(n23240) );
  MUX2S U17486 ( .A(gray_img[934]), .B(gray_img[806]), .S(n28804), .O(n25762)
         );
  MUX2S U17487 ( .A(gray_img[390]), .B(gray_img[262]), .S(n23360), .O(n18135)
         );
  NR2 U17488 ( .I1(n29680), .I2(n18134), .O(n30128) );
  MUX2S U17489 ( .A(gray_img[910]), .B(gray_img[782]), .S(n29629), .O(n29644)
         );
  ND2S U17490 ( .I1(n20907), .I2(n25374), .O(n30103) );
  MUX2S U17491 ( .A(gray_img[694]), .B(gray_img[566]), .S(n28215), .O(n28181)
         );
  ND2S U17492 ( .I1(n20952), .I2(n25374), .O(n28248) );
  MUX2S U17493 ( .A(gray_img[550]), .B(gray_img[678]), .S(n28679), .O(n28644)
         );
  ND2S U17494 ( .I1(n20935), .I2(n25374), .O(n28707) );
  OR2 U17495 ( .I1(n29680), .I2(n28642), .O(n28712) );
  MUX2S U17496 ( .A(gray_img[534]), .B(gray_img[662]), .S(n29081), .O(n29096)
         );
  ND2S U17497 ( .I1(n21006), .I2(n25374), .O(n29374) );
  MUX2S U17498 ( .A(gray_img[654]), .B(gray_img[526]), .S(n29930), .O(n29945)
         );
  MUX2S U17499 ( .A(gray_img[158]), .B(gray_img[30]), .S(n27877), .O(n27888)
         );
  ND2S U17500 ( .I1(n20964), .I2(n25374), .O(n30081) );
  NR2 U17501 ( .I1(n29680), .I2(n27887), .O(n30087) );
  MUX2S U17502 ( .A(gray_img[318]), .B(gray_img[446]), .S(n26514), .O(n26528)
         );
  ND2S U17503 ( .I1(n25087), .I2(n25374), .O(n27845) );
  MUX2S U17504 ( .A(gray_img[294]), .B(gray_img[422]), .S(n27288), .O(n27303)
         );
  MUX2S U17505 ( .A(gray_img[62]), .B(gray_img[190]), .S(n27735), .O(n27750)
         );
  MUX2S U17506 ( .A(gray_img[166]), .B(gray_img[38]), .S(n26969), .O(n26984)
         );
  ND2S U17507 ( .I1(n25275), .I2(n25374), .O(n27371) );
  MUX2S U17508 ( .A(gray_img[1998]), .B(gray_img[1870]), .S(n23582), .O(n25637) );
  ND2S U17509 ( .I1(n23584), .I2(n25374), .O(n25751) );
  NR2 U17510 ( .I1(n29680), .I2(n23581), .O(n25758) );
  MUX2S U17511 ( .A(gray_img[926]), .B(gray_img[798]), .S(n29299), .O(n29314)
         );
  ND2S U17512 ( .I1(n20940), .I2(n25374), .O(n23195) );
  NR2 U17513 ( .I1(n29680), .I2(n23161), .O(n23194) );
  MUX2S U17514 ( .A(gray_img[1966]), .B(gray_img[1838]), .S(n30018), .O(n26693) );
  ND2S U17515 ( .I1(n20958), .I2(n25374), .O(n30021) );
  MUX2S U17516 ( .A(gray_img[1950]), .B(gray_img[1822]), .S(n29517), .O(n29530) );
  MUX2S U17517 ( .A(gray_img[1934]), .B(gray_img[1806]), .S(n29415), .O(n29426) );
  ND2S U17518 ( .I1(n25219), .I2(n25374), .O(n30092) );
  MUX2S U17519 ( .A(gray_img[1790]), .B(gray_img[1662]), .S(n26009), .O(n26024) );
  ND2S U17520 ( .I1(n25082), .I2(n25374), .O(n26073) );
  MUX2S U17521 ( .A(gray_img[1646]), .B(gray_img[1774]), .S(n25805), .O(n25820) );
  ND2S U17522 ( .I1(n21077), .I2(n25374), .O(n25929) );
  ND2S U17523 ( .I1(n20895), .I2(n25374), .O(n25605) );
  MUX2S U17524 ( .A(gray_img[1614]), .B(gray_img[1742]), .S(n25679), .O(n25694) );
  ND2S U17525 ( .I1(n25025), .I2(n25374), .O(n25744) );
  MUX2S U17526 ( .A(gray_img[1718]), .B(gray_img[1590]), .S(n29222), .O(n29233) );
  ND2S U17527 ( .I1(n21083), .I2(n25374), .O(n29266) );
  MUX2S U17528 ( .A(gray_img[1710]), .B(gray_img[1582]), .S(n29121), .O(n29136) );
  MUX2S U17529 ( .A(gray_img[1686]), .B(gray_img[1558]), .S(n29577), .O(n26570) );
  ND2S U17530 ( .I1(n25096), .I2(n25374), .O(n29580) );
  MUX2S U17531 ( .A(gray_img[1678]), .B(gray_img[1550]), .S(n26601), .O(n26616) );
  ND2S U17532 ( .I1(n25104), .I2(n25374), .O(n29481) );
  MUX2S U17533 ( .A(gray_img[1398]), .B(gray_img[1526]), .S(n28134), .O(n27929) );
  ND2S U17534 ( .I1(n25284), .I2(n25374), .O(n28137) );
  INV1S U17535 ( .I(n27927), .O(n27928) );
  OR2 U17536 ( .I1(n29680), .I2(n27927), .O(n28142) );
  MUX2S U17537 ( .A(gray_img[1518]), .B(gray_img[1390]), .S(n28003), .O(n28018) );
  MUX2S U17538 ( .A(gray_img[1374]), .B(gray_img[1502]), .S(n28385), .O(n28400) );
  ND2S U17539 ( .I1(n23538), .I2(n25374), .O(n28581) );
  NR2 U17540 ( .I1(n29680), .I2(n23535), .O(n28588) );
  MUX2S U17541 ( .A(gray_img[1462]), .B(gray_img[1334]), .S(n18084), .O(n18093) );
  ND2S U17542 ( .I1(n18096), .I2(n25374), .O(n29344) );
  MUX2S U17543 ( .A(gray_img[1454]), .B(gray_img[1326]), .S(n28975), .O(n28988) );
  ND2S U17544 ( .I1(n21059), .I2(n25374), .O(n29033) );
  MUX2S U17545 ( .A(gray_img[1302]), .B(gray_img[1430]), .S(n29773), .O(n29788) );
  ND2S U17546 ( .I1(n25309), .I2(n25374), .O(n29898) );
  MUX2S U17547 ( .A(gray_img[1294]), .B(gray_img[1422]), .S(n29991), .O(n29681) );
  ND2S U17548 ( .I1(n20946), .I2(n25374), .O(n29994) );
  NR2 U17549 ( .I1(n29680), .I2(n29679), .O(n29993) );
  INV1S U17550 ( .I(n29678), .O(n29679) );
  OR2 U17551 ( .I1(n29680), .I2(n29678), .O(n29999) );
  ND2S U17552 ( .I1(n20924), .I2(n25374), .O(n23493) );
  INV1S U17553 ( .I(n23333), .O(n23334) );
  MUX2S U17554 ( .A(gray_img[1278]), .B(gray_img[1150]), .S(n23490), .O(n23350) );
  MUX2S U17555 ( .A(gray_img[1134]), .B(gray_img[1262]), .S(n28056), .O(n28069) );
  MUX2S U17556 ( .A(gray_img[1246]), .B(gray_img[1118]), .S(n28315), .O(n28330) );
  MUX2S U17557 ( .A(gray_img[1222]), .B(gray_img[1094]), .S(n28669), .O(n28518) );
  ND2S U17558 ( .I1(n25196), .I2(n25374), .O(n28672) );
  MUX2S U17559 ( .A(gray_img[1214]), .B(gray_img[1086]), .S(n28879), .O(n28894) );
  ND2S U17560 ( .I1(n20889), .I2(n25374), .O(n29044) );
  MUX2S U17561 ( .A(gray_img[1198]), .B(gray_img[1070]), .S(n29041), .O(n26140) );
  ND2S U17562 ( .I1(n25138), .I2(n25374), .O(n29881) );
  MUX2S U17563 ( .A(gray_img[1174]), .B(gray_img[1046]), .S(n29853), .O(n29823) );
  MUX2S U17564 ( .A(gray_img[1158]), .B(gray_img[1030]), .S(n29731), .O(n26651) );
  ND2S U17565 ( .I1(n25110), .I2(n25374), .O(n29740) );
  MUX2S U17566 ( .A(gray_img[886]), .B(gray_img[1014]), .S(n26401), .O(n26416)
         );
  ND2S U17567 ( .I1(n21012), .I2(n25374), .O(n26466) );
  MUX2S U17568 ( .A(gray_img[1006]), .B(gray_img[878]), .S(n26256), .O(n26271)
         );
  ND2S U17569 ( .I1(n23090), .I2(n25374), .O(n25151) );
  NR2 U17570 ( .I1(n29680), .I2(n23087), .O(n23121) );
  INV1S U17571 ( .I(n23086), .O(n23087) );
  MUX2S U17572 ( .A(gray_img[862]), .B(gray_img[990]), .S(n23088), .O(n23115)
         );
  OR2 U17573 ( .I1(n29680), .I2(n23086), .O(n23126) );
  NR2 U17574 ( .I1(n29680), .I2(n23004), .O(n27226) );
  ND2 U17575 ( .I1(n15869), .I2(n23004), .O(n27230) );
  MUX2S U17576 ( .A(gray_img[758]), .B(gray_img[630]), .S(n26360), .O(n26370)
         );
  ND2S U17577 ( .I1(n20970), .I2(n25374), .O(n26483) );
  NR2 U17578 ( .I1(n29680), .I2(n26369), .O(n26489) );
  MUX2S U17579 ( .A(n15904), .B(n26322), .S(gray_img[310]), .O(n26206) );
  ND2 U17580 ( .I1(n26207), .I2(n15869), .O(n26331) );
  MUX2S U17581 ( .A(gray_img[598]), .B(gray_img[726]), .S(n27038), .O(n27053)
         );
  ND2S U17582 ( .I1(n20901), .I2(n25374), .O(n27114) );
  ND2S U17583 ( .I1(n25163), .I2(n25374), .O(n27252) );
  MUX2S U17584 ( .A(gray_img[718]), .B(gray_img[590]), .S(n27244), .O(n27170)
         );
  INV1S U17585 ( .I(n27252), .O(n27254) );
  MUX2S U17586 ( .A(gray_img[510]), .B(gray_img[382]), .S(n27623), .O(n27636)
         );
  MUX2S U17587 ( .A(gray_img[366]), .B(gray_img[494]), .S(n27476), .O(n27491)
         );
  ND2S U17588 ( .I1(n25247), .I2(n25374), .O(n27356) );
  MUX2S U17589 ( .A(gray_img[478]), .B(gray_img[350]), .S(n27353), .O(n26798)
         );
  MUX2S U17590 ( .A(gray_img[462]), .B(gray_img[334]), .S(n23410), .O(n26867)
         );
  NR2 U17591 ( .I1(n29680), .I2(n23409), .O(n26939) );
  MUX2S U17592 ( .A(gray_img[246]), .B(gray_img[118]), .S(n27586), .O(n27598)
         );
  MUX2S U17593 ( .A(gray_img[238]), .B(gray_img[110]), .S(n27421), .O(n27436)
         );
  ND2S U17594 ( .I1(n25127), .I2(n25374), .O(n27550) );
  MUX2S U17595 ( .A(gray_img[214]), .B(gray_img[86]), .S(n23483), .O(n26731)
         );
  MUX2S U17596 ( .A(gray_img[198]), .B(gray_img[70]), .S(n23624), .O(n23632)
         );
  ND2S U17597 ( .I1(n23626), .I2(n25374), .O(n26924) );
  MUX2S U17598 ( .A(gray_img[1886]), .B(gray_img[2014]), .S(n23276), .O(n25482) );
  ND2S U17599 ( .I1(n23288), .I2(n25374), .O(n25612) );
  ND2S U17600 ( .I1(n19915), .I2(n16048), .O(n20634) );
  ND2S U17601 ( .I1(n19865), .I2(n16048), .O(n20623) );
  ND2S U17602 ( .I1(n19874), .I2(n16048), .O(n20483) );
  ND2S U17603 ( .I1(n19714), .I2(n16048), .O(n20260) );
  ND2S U17604 ( .I1(n19721), .I2(n16048), .O(n20499) );
  ND2S U17605 ( .I1(n19904), .I2(n16048), .O(n20628) );
  ND2S U17606 ( .I1(n23453), .I2(n25374), .O(n30114) );
  MUX2S U17607 ( .A(gray_img[6]), .B(gray_img[134]), .S(n23444), .O(n23473) );
  NR2 U17608 ( .I1(n29680), .I2(n23451), .O(n30120) );
  INV1S U17609 ( .I(n23450), .O(n23451) );
  INV1S U17610 ( .I(cnt_dyn[1]), .O(n30349) );
  MUX2S U17611 ( .A(n30050), .B(n20743), .S(gray_img[1088]), .O(n19134) );
  MOAI1S U17612 ( .A1(n17640), .A2(n26174), .B1(n17758), .B2(gray_img[871]), 
        .O(n16170) );
  INV2 U17613 ( .I(n17221), .O(n17079) );
  INV2 U17614 ( .I(n16165), .O(n17640) );
  INV3 U17615 ( .I(n17704), .O(n17767) );
  OR2S U17616 ( .I1(n16198), .I2(n16209), .O(n16003) );
  OR2S U17617 ( .I1(n16208), .I2(n16174), .O(n16461) );
  OR2S U17618 ( .I1(n16168), .I2(n16173), .O(n15940) );
  INV1S U17619 ( .I(n23713), .O(n23714) );
  NR2 U17620 ( .I1(n24232), .I2(n24225), .O(n24235) );
  ND2S U17621 ( .I1(n24445), .I2(n24447), .O(n24231) );
  OAI12HS U17622 ( .B1(n24229), .B2(n24228), .A1(n24227), .O(n24234) );
  NR2 U17623 ( .I1(n24148), .I2(n24142), .O(n24151) );
  NR2 U17624 ( .I1(n24605), .I2(n23956), .O(n23706) );
  NR2 U17625 ( .I1(n23653), .I2(n23687), .O(n23665) );
  NR2 U17626 ( .I1(n23655), .I2(n23687), .O(n23662) );
  OAI12HS U17627 ( .B1(n24128), .B2(n24127), .A1(n24126), .O(n24133) );
  ND2S U17628 ( .I1(n16787), .I2(cnt_cro_3b3[0]), .O(n16790) );
  AO222S U17629 ( .A1(template_reg[38]), .A2(n17581), .B1(template_reg[46]), 
        .B2(n17580), .C1(n17579), .C2(template_reg[30]), .O(n16787) );
  ND2S U17630 ( .I1(n16975), .I2(cnt_cro_3b3[0]), .O(n16978) );
  AO222S U17631 ( .A1(template_reg[37]), .A2(n17581), .B1(template_reg[45]), 
        .B2(n17580), .C1(n17579), .C2(template_reg[29]), .O(n16975) );
  BUF2 U17632 ( .I(n16182), .O(n17785) );
  INV2 U17633 ( .I(n17709), .O(n17745) );
  INV2 U17634 ( .I(n16265), .O(n17780) );
  BUF2 U17635 ( .I(n16189), .O(n17778) );
  ND2P U17636 ( .I1(n16172), .I2(n16171), .O(n17760) );
  BUF2 U17637 ( .I(n16183), .O(n17787) );
  INV2 U17638 ( .I(n16265), .O(n17591) );
  BUF2 U17639 ( .I(n16206), .O(n17797) );
  BUF2 U17640 ( .I(n16167), .O(n17759) );
  BUF2 U17641 ( .I(n16166), .O(n17758) );
  INV2 U17642 ( .I(n17221), .O(n17770) );
  ND2S U17643 ( .I1(n16070), .I2(n30375), .O(n16103) );
  OAI12HS U17644 ( .B1(n23860), .B2(n23859), .A1(n23858), .O(n23891) );
  ND2S U17645 ( .I1(n23848), .I2(n23857), .O(n23859) );
  AOI12HS U17646 ( .B1(n23887), .B2(n23886), .A1(n23885), .O(n23888) );
  ND2S U17647 ( .I1(n23878), .I2(n23887), .O(n23889) );
  AOI12HS U17648 ( .B1(n23875), .B2(n23874), .A1(n23873), .O(n23890) );
  ND2S U17649 ( .I1(n24240), .I2(n24518), .O(n24242) );
  AN2 U17650 ( .I1(n24342), .I2(n24602), .O(n23956) );
  MAO222S U17651 ( .A1(n28752), .B1(gray_img[284]), .C1(n28751), .O(n28756) );
  MAO222S U17652 ( .A1(n28750), .B1(gray_img[283]), .C1(n28749), .O(n28751) );
  ND3S U17653 ( .I1(n16047), .I2(n19127), .I3(n16009), .O(n18476) );
  OR3S U17654 ( .I1(medfilt_state_d1[1]), .I2(medfilt_state_d1[0]), .I3(
        medfilt_state_d1[2]), .O(n16008) );
  OR2S U17655 ( .I1(n23842), .I2(n23905), .O(n24340) );
  ND3S U17656 ( .I1(n23811), .I2(n23810), .I3(n23809), .O(n24286) );
  INV1S U17657 ( .I(n24286), .O(n24550) );
  OR2S U17658 ( .I1(n23802), .I2(n23905), .O(n23719) );
  INV1S U17659 ( .I(n24277), .O(n24545) );
  OR2S U17660 ( .I1(n23831), .I2(n23905), .O(n23724) );
  ND3S U17661 ( .I1(n23835), .I2(n23834), .I3(n23833), .O(n24320) );
  ND3S U17662 ( .I1(n23830), .I2(n23829), .I3(n23828), .O(n24312) );
  NR2 U17663 ( .I1(n24122), .I2(n24121), .O(n24196) );
  NR2 U17664 ( .I1(n23674), .I2(n23673), .O(n24268) );
  OR2S U17665 ( .I1(n23837), .I2(n23905), .O(n23730) );
  INV2 U17666 ( .I(n17166), .O(n17957) );
  AO222S U17667 ( .A1(template_reg[12]), .A2(n17581), .B1(template_reg[4]), 
        .B2(n17579), .C1(n17580), .C2(template_reg[20]), .O(n16596) );
  ND3S U17668 ( .I1(n16594), .I2(n16593), .I3(n16592), .O(n16595) );
  AO222S U17669 ( .A1(template_reg[34]), .A2(n17581), .B1(template_reg[42]), 
        .B2(n17580), .C1(n17579), .C2(template_reg[26]), .O(n16091) );
  BUF2 U17670 ( .I(n16153), .O(n17750) );
  NR2 U17671 ( .I1(n24060), .I2(n24053), .O(n24063) );
  OAI12HS U17672 ( .B1(n24732), .B2(n24731), .A1(n24730), .O(n24734) );
  NR2 U17673 ( .I1(n23949), .I2(n24430), .O(n23938) );
  NR2 U17674 ( .I1(n23891), .I2(n24427), .O(n23946) );
  ND3S U17675 ( .I1(n23841), .I2(n23840), .I3(n23839), .O(n24273) );
  ND3S U17676 ( .I1(n23817), .I2(n23816), .I3(n23815), .O(n24296) );
  OAI12HP U17677 ( .B1(n23801), .B2(n23800), .A1(n23799), .O(n24427) );
  ND2 U17678 ( .I1(n23798), .I2(n23789), .O(n23800) );
  AOI12HS U17679 ( .B1(n23766), .B2(n23765), .A1(n23764), .O(n23801) );
  NR2P U17680 ( .I1(n23645), .I2(n23644), .O(n23914) );
  ND2S U17681 ( .I1(n24794), .I2(n24793), .O(n24707) );
  OA12S U17682 ( .B1(n28374), .B2(n22797), .A1(n22295), .O(n22298) );
  MAO222S U17683 ( .A1(gray_img[1497]), .B1(gray_img[1496]), .C1(n28360), .O(
        n28361) );
  MAO222S U17684 ( .A1(n28306), .B1(gray_img[1235]), .C1(n28305), .O(n28307)
         );
  MAO222S U17685 ( .A1(n28304), .B1(gray_img[1234]), .C1(n28303), .O(n28305)
         );
  MAO222S U17686 ( .A1(n28485), .B1(gray_img[1227]), .C1(n28484), .O(n28486)
         );
  MAO222S U17687 ( .A1(n28483), .B1(gray_img[1226]), .C1(n28482), .O(n28484)
         );
  MAO222S U17688 ( .A1(gray_img[1876]), .B1(n23266), .C1(n23265), .O(n23267)
         );
  MAO222S U17689 ( .A1(n23264), .B1(gray_img[1875]), .C1(n23263), .O(n23265)
         );
  NR2 U17690 ( .I1(cnt_dyn_d1[3]), .I2(n18455), .O(n16052) );
  AO12S U17691 ( .B1(n24208), .B2(n24207), .A1(n24206), .O(n24486) );
  OR2S U17692 ( .I1(n24637), .I2(n24693), .O(n24643) );
  OR2S U17693 ( .I1(n24638), .I2(n24695), .O(n24642) );
  OA112 U17694 ( .C1(n24620), .C2(n24554), .A1(n24553), .B1(n24552), .O(n24752) );
  ND2S U17695 ( .I1(n24761), .I2(n24277), .O(n24279) );
  OA112 U17696 ( .C1(n24620), .C2(n24540), .A1(n24539), .B1(n24538), .O(n24747) );
  OR2S U17697 ( .I1(n23946), .I2(n23939), .O(n23967) );
  OR2S U17698 ( .I1(n23938), .I2(n23937), .O(n23966) );
  OAI12HS U17699 ( .B1(n23781), .B2(n24270), .A1(n23771), .O(n24609) );
  ND2S U17700 ( .I1(n24639), .I2(n24170), .O(n24198) );
  AO222S U17701 ( .A1(template_reg[15]), .A2(n17581), .B1(template_reg[7]), 
        .B2(n17579), .C1(n17580), .C2(template_reg[23]), .O(n16602) );
  FA1S U17702 ( .A(cro_mac[12]), .B(n17975), .CI(n17974), .CO(n17983), .S(
        n17978) );
  AO222S U17703 ( .A1(template_reg[11]), .A2(n17581), .B1(template_reg[3]), 
        .B2(n17579), .C1(n17580), .C2(template_reg[19]), .O(n16402) );
  ND3S U17704 ( .I1(n17361), .I2(n17360), .I3(n17359), .O(n17362) );
  ND3S U17705 ( .I1(n17742), .I2(n17741), .I3(n17740), .O(n17820) );
  NR2 U17706 ( .I1(n16391), .I2(n16390), .O(n17817) );
  NR2 U17707 ( .I1(n16391), .I2(n16339), .O(n17819) );
  NR2 U17708 ( .I1(n16340), .I2(n16390), .O(n17688) );
  AO222S U17709 ( .A1(template_reg[32]), .A2(n17581), .B1(template_reg[40]), 
        .B2(n17580), .C1(n17579), .C2(template_reg[24]), .O(n17582) );
  NR2 U17710 ( .I1(cnt_cro_3b3[1]), .I2(n24940), .O(n17580) );
  OR2 U17711 ( .I1(n24429), .I2(n24761), .O(n24434) );
  OR2S U17712 ( .I1(n23995), .I2(n24041), .O(n23999) );
  MAOI1S U17713 ( .A1(n23689), .A2(mem_data_out_reg_shift_1[16]), .B1(n23688), 
        .B2(n23687), .O(n23908) );
  NR2P U17714 ( .I1(n23895), .I2(n23896), .O(n24429) );
  ND2 U17715 ( .I1(n24198), .I2(n24197), .O(n24188) );
  INV1S U17716 ( .I(n24205), .O(n24160) );
  NR2P U17717 ( .I1(n24639), .I2(n24382), .O(n24208) );
  OA12S U17718 ( .B1(n24335), .B2(n24334), .A1(n24333), .O(n24336) );
  OR2S U17719 ( .I1(n24335), .I2(n24332), .O(n24337) );
  OAI12HS U17720 ( .B1(n23781), .B2(n24265), .A1(n23751), .O(n24556) );
  INV1S U17721 ( .I(n24296), .O(n24560) );
  NR2 U17722 ( .I1(n24427), .I2(n24429), .O(n24610) );
  INV1S U17723 ( .I(n22658), .O(n22619) );
  ND2S U17724 ( .I1(n30299), .I2(n30330), .O(n21131) );
  INV1S U17725 ( .I(gray_img[57]), .O(n27709) );
  OR2S U17726 ( .I1(n21151), .I2(n21158), .O(n22803) );
  ND2S U17727 ( .I1(n30451), .I2(cnt_bdyn[3]), .O(n21144) );
  ND2S U17728 ( .I1(n30132), .I2(n30365), .O(n21156) );
  ND3S U17729 ( .I1(n21745), .I2(n21744), .I3(n21743), .O(n21746) );
  OR2S U17730 ( .I1(n21146), .I2(n21138), .O(n22383) );
  ND2S U17731 ( .I1(cnt_bdyn[3]), .I2(n30298), .O(n21159) );
  ND2S U17732 ( .I1(cnt_bdyn[2]), .I2(n30132), .O(n21158) );
  ND2S U17733 ( .I1(n30302), .I2(n30365), .O(n21157) );
  ND2S U17734 ( .I1(cnt_bdyn[3]), .I2(n30424), .O(n21154) );
  MAO222 U17735 ( .A1(n28795), .B1(n28793), .C1(n28767), .O(n28768) );
  MAO222 U17736 ( .A1(n28800), .B1(n28798), .C1(n28766), .O(n28767) );
  MAO222 U17737 ( .A1(n28817), .B1(n28843), .C1(n28846), .O(n28766) );
  MAO222 U17738 ( .A1(n28226), .B1(n28230), .C1(n26126), .O(n26127) );
  MAO222S U17739 ( .A1(n28231), .B1(n28235), .C1(n26125), .O(n26126) );
  MAO222S U17740 ( .A1(n28734), .B1(n28245), .C1(n28241), .O(n26125) );
  MAO222S U17741 ( .A1(n25963), .B1(gray_img[1908]), .C1(n25962), .O(n25964)
         );
  MAO222S U17742 ( .A1(n25961), .B1(gray_img[1907]), .C1(n25960), .O(n25962)
         );
  MAO222S U17743 ( .A1(n25959), .B1(gray_img[1906]), .C1(n25958), .O(n25960)
         );
  AO22S U17744 ( .A1(n26060), .A2(n26062), .B1(n25973), .B2(n15979), .O(n15968) );
  OR2S U17745 ( .I1(n26060), .I2(n26062), .O(n15979) );
  MAO222 U17746 ( .A1(n26067), .B1(n26065), .C1(n25972), .O(n25973) );
  MAO222 U17747 ( .A1(n26072), .B1(n26070), .C1(n25971), .O(n25972) );
  MAO222 U17748 ( .A1(n25922), .B1(n25920), .C1(n25863), .O(n25864) );
  MAO222 U17749 ( .A1(n25927), .B1(n25925), .C1(n25862), .O(n25863) );
  MAO222 U17750 ( .A1(n26095), .B1(n25939), .C1(n25941), .O(n25862) );
  MAO222S U17751 ( .A1(n23226), .B1(gray_img[804]), .C1(n23225), .O(n23227) );
  MAO222S U17752 ( .A1(n23224), .B1(gray_img[803]), .C1(n23223), .O(n23225) );
  MAO222 U17753 ( .A1(n28695), .B1(n28699), .C1(n23234), .O(n23235) );
  MAO222S U17754 ( .A1(n28700), .B1(n28704), .C1(n23233), .O(n23234) );
  MAO222S U17755 ( .A1(n28813), .B1(n23246), .C1(n23241), .O(n23233) );
  MAO222S U17756 ( .A1(n18107), .B1(gray_img[268]), .C1(n18106), .O(n18108) );
  MAO222S U17757 ( .A1(n18105), .B1(gray_img[267]), .C1(n18104), .O(n18106) );
  MAO222 U17758 ( .A1(n30055), .B1(n30053), .C1(n18128), .O(n18129) );
  MAO222S U17759 ( .A1(n30062), .B1(n30060), .C1(n18127), .O(n18128) );
  MAO222S U17760 ( .A1(n29622), .B1(gray_img[772]), .C1(n29621), .O(n29623) );
  MAO222S U17761 ( .A1(n29620), .B1(gray_img[771]), .C1(n29619), .O(n29621) );
  MAO222 U17762 ( .A1(n29985), .B1(n29983), .C1(n29631), .O(n29632) );
  MAO222 U17763 ( .A1(n29990), .B1(n29988), .C1(n29630), .O(n29631) );
  MAO222S U17764 ( .A1(n30017), .B1(n30015), .C1(n30108), .O(n29630) );
  MAO222 U17765 ( .A1(n28191), .B1(n28195), .C1(n28172), .O(n28173) );
  MAO222 U17766 ( .A1(n28196), .B1(n28200), .C1(n28171), .O(n28172) );
  MAO222S U17767 ( .A1(n28220), .B1(n28240), .C1(n28236), .O(n28171) );
  MAO222 U17768 ( .A1(n28659), .B1(n28663), .C1(n28635), .O(n28636) );
  MAO222S U17769 ( .A1(n28664), .B1(n28668), .C1(n28634), .O(n28635) );
  MAO222S U17770 ( .A1(n28684), .B1(n28713), .C1(n28705), .O(n28634) );
  MAO222S U17771 ( .A1(n29054), .B1(gray_img[659]), .C1(n29053), .O(n29055) );
  MAO222S U17772 ( .A1(intadd_132_B_1_), .B1(gray_img[658]), .C1(n29052), .O(
        n29053) );
  MAO222S U17773 ( .A1(n29070), .B1(gray_img[668]), .C1(n29069), .O(n29075) );
  MAO222S U17774 ( .A1(n29068), .B1(gray_img[667]), .C1(n29067), .O(n29069) );
  MAO222S U17775 ( .A1(n29066), .B1(gray_img[666]), .C1(n29065), .O(n29067) );
  MAO222S U17776 ( .A1(n29334), .B1(n29332), .C1(n29083), .O(n29084) );
  MAO222 U17777 ( .A1(n29339), .B1(n29337), .C1(n29082), .O(n29083) );
  MAO222 U17778 ( .A1(n29358), .B1(n29377), .C1(n29380), .O(n29082) );
  MAO222S U17779 ( .A1(n29921), .B1(gray_img[643]), .C1(n29920), .O(n29922) );
  MAO222S U17780 ( .A1(n29919), .B1(gray_img[642]), .C1(n29918), .O(n29920) );
  MAO222S U17781 ( .A1(intadd_8_B_0_), .B1(gray_img[641]), .C1(intadd_8_CI), 
        .O(n29918) );
  MAO222 U17782 ( .A1(n29960), .B1(n29958), .C1(n29932), .O(n29933) );
  MAO222 U17783 ( .A1(n29965), .B1(n29963), .C1(n29931), .O(n29932) );
  MAO222 U17784 ( .A1(n30011), .B1(n29968), .C1(n29970), .O(n29931) );
  MAO222 U17785 ( .A1(n28834), .B1(n28832), .C1(n27879), .O(n27880) );
  MAO222 U17786 ( .A1(n28839), .B1(n28837), .C1(n27878), .O(n27879) );
  MAO222S U17787 ( .A1(n28852), .B1(n28850), .C1(n30086), .O(n27878) );
  MAO222S U17788 ( .A1(n26507), .B1(gray_img[436]), .C1(n26506), .O(n26508) );
  MAO222S U17789 ( .A1(n26505), .B1(gray_img[435]), .C1(n26504), .O(n26506) );
  MAO222S U17790 ( .A1(n26503), .B1(gray_img[434]), .C1(n26502), .O(n26504) );
  AO22S U17791 ( .A1(n27806), .A2(n27808), .B1(n26516), .B2(n15977), .O(n15978) );
  MAO222 U17792 ( .A1(n27813), .B1(n27811), .C1(n26515), .O(n26516) );
  MAO222 U17793 ( .A1(n27850), .B1(n27824), .C1(n27826), .O(n26515) );
  MAO222 U17794 ( .A1(n27269), .B1(gray_img[420]), .C1(n27268), .O(n27270) );
  MAO222S U17795 ( .A1(gray_img[291]), .B1(n27266), .C1(n27265), .O(n27267) );
  MAO222 U17796 ( .A1(n27319), .B1(n27317), .C1(n27290), .O(n27291) );
  MAO222 U17797 ( .A1(n27324), .B1(n27322), .C1(n27289), .O(n27290) );
  MAO222 U17798 ( .A1(n30075), .B1(n27327), .C1(n27329), .O(n27289) );
  MAO222 U17799 ( .A1(n27766), .B1(n27764), .C1(n27737), .O(n27738) );
  MAO222S U17800 ( .A1(n27771), .B1(n27769), .C1(n27736), .O(n27737) );
  MAO222 U17801 ( .A1(n27820), .B1(n27817), .C1(n27793), .O(n27736) );
  MAO222 U17802 ( .A1(n26949), .B1(gray_img[36]), .C1(n26948), .O(n26950) );
  MAO222S U17803 ( .A1(n26947), .B1(gray_img[35]), .C1(n26946), .O(n26948) );
  MAO222S U17804 ( .A1(n26962), .B1(gray_img[172]), .C1(n26961), .O(n26963) );
  MAO222S U17805 ( .A1(n26960), .B1(gray_img[171]), .C1(n26959), .O(n26961) );
  MAO222S U17806 ( .A1(n26958), .B1(gray_img[170]), .C1(n26957), .O(n26959) );
  MAO222 U17807 ( .A1(n27344), .B1(n27342), .C1(n26971), .O(n26972) );
  MAO222 U17808 ( .A1(n27349), .B1(n27347), .C1(n26970), .O(n26971) );
  MAO222S U17809 ( .A1(n27370), .B1(n27374), .C1(n27377), .O(n26970) );
  MAO222S U17810 ( .A1(n29280), .B1(gray_img[796]), .C1(n29279), .O(n29281) );
  MAO222S U17811 ( .A1(n29278), .B1(gray_img[795]), .C1(n29277), .O(n29279) );
  MAO222 U17812 ( .A1(n29368), .B1(n29366), .C1(n29301), .O(n29302) );
  MAO222 U17813 ( .A1(n29373), .B1(n29371), .C1(n29300), .O(n29301) );
  MAO222S U17814 ( .A1(n30037), .B1(n29384), .C1(n29386), .O(n29300) );
  MAO222S U17815 ( .A1(n23132), .B1(gray_img[1852]), .C1(n23131), .O(n23133)
         );
  MAO222S U17816 ( .A1(n23130), .B1(gray_img[1851]), .C1(n23129), .O(n23131)
         );
  MAO222S U17817 ( .A1(intadd_159_B_1_), .B1(gray_img[1850]), .C1(n23128), .O(
        n23129) );
  MAO222S U17818 ( .A1(n23144), .B1(gray_img[1844]), .C1(n23143), .O(n23145)
         );
  MAO222 U17819 ( .A1(n23168), .B1(n23172), .C1(n23153), .O(n23154) );
  MAO222 U17820 ( .A1(n23173), .B1(n23177), .C1(n23152), .O(n23153) );
  MAO222S U17821 ( .A1(n23201), .B1(n23167), .C1(n23193), .O(n23152) );
  MAO222 U17822 ( .A1(n29172), .B1(n29176), .C1(n26684), .O(n26685) );
  MAO222S U17823 ( .A1(n29177), .B1(n29181), .C1(n26683), .O(n26684) );
  MAO222S U17824 ( .A1(n29197), .B1(n30027), .C1(n29193), .O(n26683) );
  MAO222S U17825 ( .A1(n29510), .B1(gray_img[1820]), .C1(n29509), .O(n29511)
         );
  MAO222S U17826 ( .A1(n29508), .B1(gray_img[1819]), .C1(n29507), .O(n29509)
         );
  MAO222S U17827 ( .A1(n29506), .B1(gray_img[1818]), .C1(n29505), .O(n29507)
         );
  AO22S U17828 ( .A1(n29563), .A2(n29565), .B1(n29520), .B2(n15971), .O(n15953) );
  OR2S U17829 ( .I1(n29563), .I2(n29565), .O(n15971) );
  MAO222 U17830 ( .A1(n29571), .B1(n29569), .C1(n29519), .O(n29520) );
  MAO222 U17831 ( .A1(n29576), .B1(n29574), .C1(n29518), .O(n29519) );
  MAO222S U17832 ( .A1(n29389), .B1(gray_img[1922]), .C1(n29388), .O(n29390)
         );
  MAO222S U17833 ( .A1(gray_img[1921]), .B1(gray_img[1920]), .C1(n29387), .O(
        n29388) );
  MAO222S U17834 ( .A1(gray_img[1805]), .B1(n29408), .C1(n29407), .O(n29410)
         );
  MAO222 U17835 ( .A1(gray_img[1804]), .B1(n29406), .C1(n29405), .O(n29407) );
  MAO222S U17836 ( .A1(gray_img[1803]), .B1(n29404), .C1(n29403), .O(n29405)
         );
  MAO222S U17837 ( .A1(gray_img[1802]), .B1(n29402), .C1(n29401), .O(n29403)
         );
  MAO222 U17838 ( .A1(n29471), .B1(n29469), .C1(n29417), .O(n29418) );
  MAO222S U17839 ( .A1(n29476), .B1(n29474), .C1(n29416), .O(n29417) );
  MAO222S U17840 ( .A1(n29492), .B1(n29490), .C1(n30097), .O(n29416) );
  MAO222S U17841 ( .A1(n26004), .B1(gray_img[1653]), .C1(n26003), .O(n26005)
         );
  MAO222S U17842 ( .A1(n26002), .B1(gray_img[1652]), .C1(n26001), .O(n26003)
         );
  MAO222S U17843 ( .A1(n26000), .B1(gray_img[1651]), .C1(n25999), .O(n26001)
         );
  MAO222 U17844 ( .A1(n26039), .B1(n26037), .C1(n26011), .O(n26012) );
  MAO222 U17845 ( .A1(n26044), .B1(n26042), .C1(n26010), .O(n26011) );
  MAO222S U17846 ( .A1(n26079), .B1(n26076), .C1(n26052), .O(n26010) );
  MAO222S U17847 ( .A1(n25784), .B1(gray_img[1771]), .C1(n25783), .O(n25785)
         );
  MAO222S U17848 ( .A1(n25782), .B1(gray_img[1770]), .C1(n25781), .O(n25783)
         );
  MAO222S U17849 ( .A1(gray_img[1769]), .B1(gray_img[1768]), .C1(n25780), .O(
        n25781) );
  MAO222 U17850 ( .A1(n25891), .B1(n25889), .C1(n25807), .O(n25808) );
  MAO222 U17851 ( .A1(n25896), .B1(n25894), .C1(n25806), .O(n25807) );
  MAO222S U17852 ( .A1(n25935), .B1(n25932), .C1(n25907), .O(n25806) );
  MAO222 U17853 ( .A1(n25564), .B1(n25568), .C1(n25540), .O(n25541) );
  MAO222S U17854 ( .A1(n25569), .B1(n25573), .C1(n25539), .O(n25540) );
  MAO222S U17855 ( .A1(n25611), .B1(n25582), .C1(n25603), .O(n25539) );
  MAO222S U17856 ( .A1(n25658), .B1(gray_img[1739]), .C1(n25657), .O(n25659)
         );
  MAO222S U17857 ( .A1(n25656), .B1(gray_img[1738]), .C1(n25655), .O(n25657)
         );
  MAO222S U17858 ( .A1(gray_img[1737]), .B1(gray_img[1736]), .C1(n25654), .O(
        n25655) );
  MAO222 U17859 ( .A1(n25709), .B1(n25707), .C1(n25681), .O(n25682) );
  MAO222 U17860 ( .A1(n25714), .B1(n25712), .C1(n25680), .O(n25681) );
  MAO222 U17861 ( .A1(n25719), .B1(n25717), .C1(n25749), .O(n25680) );
  MAO222 U17862 ( .A1(n29252), .B1(n29250), .C1(n29224), .O(n29225) );
  MAO222 U17863 ( .A1(n29257), .B1(n29255), .C1(n29223), .O(n29224) );
  MAO222S U17864 ( .A1(n29272), .B1(n29269), .C1(n29265), .O(n29223) );
  MAO222 U17865 ( .A1(n29151), .B1(n29149), .C1(n29123), .O(n29124) );
  MAO222 U17866 ( .A1(n29156), .B1(n29154), .C1(n29122), .O(n29123) );
  MAO222S U17867 ( .A1(n29161), .B1(n29159), .C1(n29191), .O(n29122) );
  MAO222S U17868 ( .A1(n29541), .B1(n29545), .C1(n26561), .O(n26562) );
  MAO222 U17869 ( .A1(n29546), .B1(n29550), .C1(n26560), .O(n26561) );
  MAO222S U17870 ( .A1(n29586), .B1(n29555), .C1(n29551), .O(n26560) );
  MAO222S U17871 ( .A1(n26581), .B1(gray_img[1548]), .C1(n26580), .O(n26582)
         );
  MAO222S U17872 ( .A1(n26579), .B1(gray_img[1547]), .C1(n26578), .O(n26580)
         );
  MAO222S U17873 ( .A1(n26577), .B1(gray_img[1546]), .C1(n26576), .O(n26578)
         );
  MAO222 U17874 ( .A1(n29446), .B1(n29444), .C1(n26603), .O(n26604) );
  MAO222S U17875 ( .A1(n29451), .B1(n29449), .C1(n26602), .O(n26603) );
  MAO222S U17876 ( .A1(n29456), .B1(n29454), .C1(n29486), .O(n26602) );
  MAO222S U17877 ( .A1(n27900), .B1(gray_img[1405]), .C1(n27899), .O(n27901)
         );
  MAO222S U17878 ( .A1(n27898), .B1(gray_img[1404]), .C1(n27897), .O(n27899)
         );
  MAO222S U17879 ( .A1(n27896), .B1(gray_img[1403]), .C1(n27895), .O(n27897)
         );
  MAO222 U17880 ( .A1(n27944), .B1(n27948), .C1(n27920), .O(n27921) );
  MAO222 U17881 ( .A1(n27949), .B1(n27953), .C1(n27919), .O(n27920) );
  MAO222S U17882 ( .A1(n28143), .B1(n27958), .C1(n27954), .O(n27919) );
  MAO222S U17883 ( .A1(n27992), .B1(gray_img[1380]), .C1(n27991), .O(n27995)
         );
  MAO222 U17884 ( .A1(n28115), .B1(n28113), .C1(n28005), .O(n28006) );
  MAO222 U17885 ( .A1(n28120), .B1(n28118), .C1(n28004), .O(n28005) );
  MAO222S U17886 ( .A1(n28133), .B1(n28131), .C1(n28213), .O(n28004) );
  MAO222 U17887 ( .A1(n28446), .B1(n28444), .C1(n28387), .O(n28388) );
  MAO222 U17888 ( .A1(n28451), .B1(n28449), .C1(n28386), .O(n28387) );
  MAO222S U17889 ( .A1(n28464), .B1(n28462), .C1(n28606), .O(n28386) );
  MAO222S U17890 ( .A1(gray_img[1349]), .B1(n23508), .C1(n23507), .O(n23509)
         );
  MAO222S U17891 ( .A1(gray_img[1348]), .B1(n23506), .C1(n23505), .O(n23507)
         );
  MAO222S U17892 ( .A1(gray_img[1347]), .B1(n23504), .C1(n23503), .O(n23505)
         );
  MAO222S U17893 ( .A1(n28547), .B1(n28545), .C1(n23528), .O(n23529) );
  MAO222 U17894 ( .A1(n28552), .B1(n28550), .C1(n23527), .O(n23528) );
  MAO222 U17895 ( .A1(n28557), .B1(n28555), .C1(n23526), .O(n23527) );
  MAO222 U17896 ( .A1(n28584), .B1(n23543), .C1(n28587), .O(n23526) );
  AO12S U17897 ( .B1(gray_img[1333]), .B2(n18075), .A1(n18074), .O(n18079) );
  MAO222S U17898 ( .A1(gray_img[1332]), .B1(n18073), .C1(n18072), .O(n18074)
         );
  MAO222 U17899 ( .A1(n28909), .B1(n28907), .C1(n18086), .O(n18087) );
  MAO222 U17900 ( .A1(n28914), .B1(n28912), .C1(n18085), .O(n18086) );
  MAO222 U17901 ( .A1(n29349), .B1(n28917), .C1(n28919), .O(n18085) );
  MAO222S U17902 ( .A1(n28968), .B1(gray_img[1324]), .C1(n28967), .O(n28969)
         );
  MAO222S U17903 ( .A1(n28966), .B1(gray_img[1323]), .C1(n28965), .O(n28967)
         );
  AO22S U17904 ( .A1(n28996), .A2(n28998), .B1(n28978), .B2(n15965), .O(n15966) );
  OR2S U17905 ( .I1(n28996), .I2(n28998), .O(n15965) );
  MAO222 U17906 ( .A1(n29003), .B1(n29001), .C1(n28977), .O(n28978) );
  MAO222 U17907 ( .A1(n29008), .B1(n29006), .C1(n28976), .O(n28977) );
  MAO222S U17908 ( .A1(n29751), .B1(gray_img[1427]), .C1(n29750), .O(n29752)
         );
  MAO222S U17909 ( .A1(n29749), .B1(gray_img[1426]), .C1(n29748), .O(n29750)
         );
  MAO222S U17910 ( .A1(intadd_62_B_0_), .B1(gray_img[1425]), .C1(n29747), .O(
        n29748) );
  MAO222S U17911 ( .A1(n29766), .B1(gray_img[1436]), .C1(n29765), .O(n29767)
         );
  MAO222S U17912 ( .A1(n29764), .B1(gray_img[1435]), .C1(n29763), .O(n29765)
         );
  MAO222S U17913 ( .A1(n29762), .B1(gray_img[1434]), .C1(n29761), .O(n29763)
         );
  MAO222 U17914 ( .A1(n29873), .B1(n29871), .C1(n29775), .O(n29776) );
  MAO222 U17915 ( .A1(n29878), .B1(n29876), .C1(n29774), .O(n29775) );
  MAO222S U17916 ( .A1(n29903), .B1(n29891), .C1(n29893), .O(n29774) );
  MAO222 U17917 ( .A1(n29696), .B1(n29700), .C1(n29671), .O(n29672) );
  MAO222 U17918 ( .A1(n29701), .B1(n29705), .C1(n29670), .O(n29671) );
  MAO222S U17919 ( .A1(n30000), .B1(n29710), .C1(n29706), .O(n29670) );
  MAO222S U17920 ( .A1(n23305), .B1(gray_img[1268]), .C1(n23304), .O(n23306)
         );
  MAO222S U17921 ( .A1(n23303), .B1(gray_img[1267]), .C1(n23302), .O(n23304)
         );
  MAO222 U17922 ( .A1(n23345), .B1(n23349), .C1(n23326), .O(n23327) );
  MAO222S U17923 ( .A1(n23335), .B1(n23339), .C1(n23325), .O(n23326) );
  MAO222S U17924 ( .A1(n23371), .B1(n23499), .C1(n23367), .O(n23325) );
  MAO222S U17925 ( .A1(n28047), .B1(gray_img[1259]), .C1(n28046), .O(n28048)
         );
  MAO222S U17926 ( .A1(n28045), .B1(gray_img[1258]), .C1(n28044), .O(n28046)
         );
  MAO222S U17927 ( .A1(gray_img[1257]), .B1(gray_img[1256]), .C1(intadd_71_CI), 
        .O(n28044) );
  AO22S U17928 ( .A1(n28077), .A2(n28079), .B1(n28059), .B2(n15963), .O(n15955) );
  MAO222 U17929 ( .A1(n28084), .B1(n28082), .C1(n28058), .O(n28059) );
  MAO222 U17930 ( .A1(n28089), .B1(n28087), .C1(n28057), .O(n28058) );
  MAO222S U17931 ( .A1(n28415), .B1(n28413), .C1(n28317), .O(n28318) );
  MAO222 U17932 ( .A1(n28420), .B1(n28418), .C1(n28316), .O(n28317) );
  MAO222 U17933 ( .A1(n28431), .B1(n28455), .C1(n28458), .O(n28316) );
  MAO222S U17934 ( .A1(n28571), .B1(n28575), .C1(n28509), .O(n28510) );
  MAO222 U17935 ( .A1(n28576), .B1(n28580), .C1(n28508), .O(n28509) );
  MAO222S U17936 ( .A1(n28678), .B1(n28593), .C1(n28589), .O(n28508) );
  MAO222S U17937 ( .A1(n28859), .B1(gray_img[1084]), .C1(n28858), .O(n28860)
         );
  MAO222S U17938 ( .A1(n28857), .B1(gray_img[1083]), .C1(n28856), .O(n28858)
         );
  MAO222 U17939 ( .A1(n28872), .B1(gray_img[1076]), .C1(n28871), .O(n28873) );
  MAO222 U17940 ( .A1(n28870), .B1(gray_img[1075]), .C1(n28869), .O(n28871) );
  MAO222 U17941 ( .A1(n28929), .B1(n28927), .C1(n28881), .O(n28882) );
  MAO222 U17942 ( .A1(n28934), .B1(n28932), .C1(n28880), .O(n28881) );
  MAO222S U17943 ( .A1(n28949), .B1(n28946), .C1(n28942), .O(n28880) );
  MAO222S U17944 ( .A1(n23012), .B1(gray_img[1059]), .C1(n23011), .O(n23013)
         );
  MAO222S U17945 ( .A1(gray_img[1057]), .B1(gray_img[1056]), .C1(intadd_83_CI), 
        .O(n23009) );
  MAO222S U17946 ( .A1(n23026), .B1(gray_img[1068]), .C1(n23025), .O(n23027)
         );
  MAO222S U17947 ( .A1(n23024), .B1(gray_img[1067]), .C1(n23023), .O(n23025)
         );
  MAO222 U17948 ( .A1(n29027), .B1(n29031), .C1(n23035), .O(n23036) );
  MAO222 U17949 ( .A1(n23044), .B1(n23048), .C1(n23034), .O(n23035) );
  MAO222 U17950 ( .A1(n23376), .B1(n29050), .C1(n23372), .O(n23034) );
  MAO222S U17951 ( .A1(n29805), .B1(gray_img[1044]), .C1(n29804), .O(n29806)
         );
  MAO222S U17952 ( .A1(n29803), .B1(gray_img[1043]), .C1(n29802), .O(n29804)
         );
  MAO222S U17953 ( .A1(intadd_85_B_1_), .B1(gray_img[1042]), .C1(n29801), .O(
        n29802) );
  MAO222 U17954 ( .A1(n29841), .B1(n29846), .C1(n29814), .O(n29815) );
  MAO222 U17955 ( .A1(n29847), .B1(n29852), .C1(n29813), .O(n29814) );
  MAO222S U17956 ( .A1(n29858), .B1(n29888), .C1(n29879), .O(n29813) );
  MAO222S U17957 ( .A1(n29721), .B1(n29725), .C1(n26642), .O(n26643) );
  MAO222 U17958 ( .A1(n29726), .B1(n29730), .C1(n26641), .O(n26642) );
  MAO222S U17959 ( .A1(n29737), .B1(n29746), .C1(n29738), .O(n26641) );
  MAO222S U17960 ( .A1(n26396), .B1(gray_img[1021]), .C1(n26395), .O(n26397)
         );
  MAO222S U17961 ( .A1(n26394), .B1(gray_img[1020]), .C1(n26393), .O(n26395)
         );
  MAO222S U17962 ( .A1(n26392), .B1(gray_img[1019]), .C1(n26391), .O(n26393)
         );
  MAO222 U17963 ( .A1(n26431), .B1(n26429), .C1(n26403), .O(n26404) );
  MAO222 U17964 ( .A1(n26436), .B1(n26434), .C1(n26402), .O(n26403) );
  MAO222S U17965 ( .A1(n26444), .B1(n26469), .C1(n26472), .O(n26402) );
  MAO222S U17966 ( .A1(gray_img[1004]), .B1(n26232), .C1(n26231), .O(n26235)
         );
  MAO222S U17967 ( .A1(n26286), .B1(n26284), .C1(n26258), .O(n26259) );
  MAO222 U17968 ( .A1(n26291), .B1(n26289), .C1(n26257), .O(n26258) );
  MAO222 U17969 ( .A1(n27839), .B1(n26294), .C1(n26296), .O(n26257) );
  MAO222 U17970 ( .A1(n23100), .B1(n23104), .C1(n23081), .O(n23082) );
  MAO222 U17971 ( .A1(n23095), .B1(n23099), .C1(n23080), .O(n23081) );
  MAO222S U17972 ( .A1(n23127), .B1(n23094), .C1(n23120), .O(n23080) );
  MAO222S U17973 ( .A1(n27198), .B1(n27201), .C1(n22993), .O(n22995) );
  MAO222 U17974 ( .A1(n27213), .B1(n27216), .C1(n22992), .O(n22993) );
  MAO222 U17975 ( .A1(n27218), .B1(n27221), .C1(n22991), .O(n22992) );
  MAO222 U17976 ( .A1(n27229), .B1(n23299), .C1(n27225), .O(n22991) );
  MAO222S U17977 ( .A1(n26338), .B1(gray_img[636]), .C1(n26337), .O(n26339) );
  MAO222S U17978 ( .A1(n26336), .B1(gray_img[635]), .C1(n26335), .O(n26337) );
  INV1S U17979 ( .I(n26359), .O(n26362) );
  MAO222 U17980 ( .A1(n26460), .B1(n26458), .C1(n26358), .O(n26359) );
  MAO222 U17981 ( .A1(n26465), .B1(n26463), .C1(n26357), .O(n26358) );
  MAO222 U17982 ( .A1(n26488), .B1(n26476), .C1(n26478), .O(n26357) );
  MAO222S U17983 ( .A1(gray_img[612]), .B1(n26168), .C1(n26167), .O(n26169) );
  MAO222S U17984 ( .A1(gray_img[611]), .B1(n26166), .C1(n26165), .O(n26167) );
  MAO222S U17985 ( .A1(gray_img[610]), .B1(n26164), .C1(n26163), .O(n26165) );
  MAO222S U17986 ( .A1(n26162), .B1(n26161), .C1(gray_img[609]), .O(n26163) );
  MAO222S U17987 ( .A1(n26303), .B1(n26306), .C1(n26193), .O(n26196) );
  MAO222 U17988 ( .A1(n26308), .B1(n26311), .C1(n26192), .O(n26193) );
  MAO222 U17989 ( .A1(n26313), .B1(n26316), .C1(n26191), .O(n26192) );
  MAO222S U17990 ( .A1(n26321), .B1(n26330), .C1(n26318), .O(n26191) );
  MAO222S U17991 ( .A1(n27017), .B1(gray_img[723]), .C1(n27016), .O(n27018) );
  MAO222S U17992 ( .A1(n27015), .B1(gray_img[722]), .C1(n27014), .O(n27016) );
  MAO222S U17993 ( .A1(gray_img[721]), .B1(gray_img[720]), .C1(intadd_105_CI), 
        .O(n27014) );
  MAO222 U17994 ( .A1(n27097), .B1(n27095), .C1(n27040), .O(n27041) );
  MAO222S U17995 ( .A1(n27102), .B1(n27100), .C1(n27039), .O(n27040) );
  MAO222S U17996 ( .A1(n27152), .B1(gray_img[588]), .C1(n27151), .O(n27153) );
  MAO222S U17997 ( .A1(n27150), .B1(gray_img[587]), .C1(n27149), .O(n27151) );
  MAO222 U17998 ( .A1(n27231), .B1(n27235), .C1(n27161), .O(n27162) );
  MAO222 U17999 ( .A1(n27236), .B1(n27240), .C1(n27160), .O(n27161) );
  MAO222S U18000 ( .A1(n27258), .B1(n27249), .C1(n27250), .O(n27160) );
  MAO222S U18001 ( .A1(n27616), .B1(gray_img[380]), .C1(n27615), .O(n27617) );
  MAO222S U18002 ( .A1(n27614), .B1(gray_img[379]), .C1(n27613), .O(n27615) );
  AO22S U18003 ( .A1(n27644), .A2(n27646), .B1(n27626), .B2(n15961), .O(n15957) );
  OR2S U18004 ( .I1(n27644), .I2(n27646), .O(n15961) );
  MAO222 U18005 ( .A1(n27651), .B1(n27649), .C1(n27625), .O(n27626) );
  MAO222 U18006 ( .A1(n27656), .B1(n27654), .C1(n27624), .O(n27625) );
  MAO222S U18007 ( .A1(n27457), .B1(gray_img[492]), .C1(n27456), .O(n27458) );
  MAO222S U18008 ( .A1(n27455), .B1(gray_img[491]), .C1(n27454), .O(n27456) );
  MAO222S U18009 ( .A1(n27453), .B1(gray_img[490]), .C1(n27452), .O(n27454) );
  MAO222 U18010 ( .A1(n27506), .B1(n27504), .C1(n27478), .O(n27479) );
  MAO222S U18011 ( .A1(n27511), .B1(n27509), .C1(n27477), .O(n27478) );
  MAO222S U18012 ( .A1(n27517), .B1(n27515), .C1(n27784), .O(n27477) );
  MAO222S U18013 ( .A1(gray_img[469]), .B1(n26770), .C1(n26769), .O(n26771) );
  MAO222S U18014 ( .A1(gray_img[468]), .B1(n26768), .C1(n26767), .O(n26769) );
  MAO222 U18015 ( .A1(n26813), .B1(n26817), .C1(n26789), .O(n26790) );
  MAO222S U18016 ( .A1(n26818), .B1(n26822), .C1(n26788), .O(n26789) );
  MAO222S U18017 ( .A1(n26827), .B1(n27362), .C1(n26823), .O(n26788) );
  MAO222S U18018 ( .A1(n23394), .B1(gray_img[332]), .C1(n23393), .O(n23395) );
  MAO222S U18019 ( .A1(n23392), .B1(gray_img[331]), .C1(n23391), .O(n23393) );
  MAO222 U18020 ( .A1(n26918), .B1(n26916), .C1(n23403), .O(n23404) );
  MAO222 U18021 ( .A1(n26923), .B1(n26921), .C1(n23402), .O(n23403) );
  MAO222S U18022 ( .A1(n26935), .B1(n23417), .C1(n26938), .O(n23402) );
  MAO222S U18023 ( .A1(n27574), .B1(gray_img[116]), .C1(n27573), .O(n27575) );
  MAO222S U18024 ( .A1(n27572), .B1(gray_img[115]), .C1(n27571), .O(n27573) );
  MAO222 U18025 ( .A1(n27674), .B1(n27672), .C1(n27583), .O(n27585) );
  MAO222 U18026 ( .A1(n27679), .B1(n27677), .C1(n27582), .O(n27583) );
  MAO222 U18027 ( .A1(n27684), .B1(n27682), .C1(n27581), .O(n27582) );
  MAO222 U18028 ( .A1(n27697), .B1(n27695), .C1(n27707), .O(n27581) );
  AO12S U18029 ( .B1(gray_img[109]), .B2(n27400), .A1(n27399), .O(n27404) );
  MAO222S U18030 ( .A1(gray_img[108]), .B1(n27398), .C1(n27397), .O(n27399) );
  MAO222S U18031 ( .A1(n27396), .B1(gray_img[107]), .C1(n27395), .O(n27397) );
  MAO222 U18032 ( .A1(n27532), .B1(n27530), .C1(n27423), .O(n27424) );
  MAO222 U18033 ( .A1(n27537), .B1(n27535), .C1(n27422), .O(n27423) );
  MAO222 U18034 ( .A1(n27555), .B1(n27540), .C1(n27542), .O(n27422) );
  MAO222S U18035 ( .A1(n16031), .B1(gray_img[84]), .C1(n16030), .O(n16032) );
  MAO222S U18036 ( .A1(n16029), .B1(gray_img[83]), .C1(n16028), .O(n16030) );
  AO22S U18037 ( .A1(n16060), .A2(n16046), .B1(n16042), .B2(n16041), .O(n15959) );
  MAO222 U18038 ( .A1(n16063), .B1(n16068), .C1(n16040), .O(n16042) );
  MAO222 U18039 ( .A1(n26898), .B1(n26896), .C1(n23617), .O(n23618) );
  MAO222 U18040 ( .A1(n26903), .B1(n26901), .C1(n23616), .O(n23617) );
  MAO222 U18041 ( .A1(n26927), .B1(n23631), .C1(n26930), .O(n23616) );
  MAO222 U18042 ( .A1(n23253), .B1(gray_img[2012]), .C1(n23252), .O(n23254) );
  MAO222S U18043 ( .A1(n23251), .B1(gray_img[2011]), .C1(n23250), .O(n23252)
         );
  MAO222S U18044 ( .A1(n23249), .B1(gray_img[2010]), .C1(n23248), .O(n23250)
         );
  MAO222S U18045 ( .A1(n25597), .B1(n25595), .C1(n23278), .O(n23279) );
  MAO222 U18046 ( .A1(n25602), .B1(n25600), .C1(n23277), .O(n23278) );
  MAO222 U18047 ( .A1(n23293), .B1(n25615), .C1(n25618), .O(n23277) );
  ND2S U18048 ( .I1(medfilt_cnt2_d1[0]), .I2(medfilt_cnt2_d1[3]), .O(n18576)
         );
  ND2S U18049 ( .I1(cnt_bdyn_d1[0]), .I2(cnt_bdyn_d1[3]), .O(n18578) );
  ND2S U18050 ( .I1(medfilt_cnt2_d1[3]), .I2(n18469), .O(n18566) );
  ND2S U18051 ( .I1(cnt_bdyn_d1[3]), .I2(n18470), .O(n18567) );
  ND2S U18052 ( .I1(medfilt_cnt2_d1[1]), .I2(medfilt_cnt2_d1[2]), .O(n18577)
         );
  ND2S U18053 ( .I1(cnt_bdyn_d1[1]), .I2(cnt_bdyn_d1[2]), .O(n18579) );
  ND2S U18054 ( .I1(medfilt_cnt2_d1[2]), .I2(n18094), .O(n18532) );
  ND2S U18055 ( .I1(cnt_bdyn_d1[2]), .I2(n18095), .O(n18533) );
  ND2S U18056 ( .I1(medfilt_cnt_d1[1]), .I2(medfilt_cnt_d1[2]), .O(n18820) );
  ND2S U18057 ( .I1(cnt_dyn_d1[1]), .I2(cnt_dyn_d1[2]), .O(n18822) );
  ND2S U18058 ( .I1(medfilt_cnt_d1[1]), .I2(n18136), .O(n24972) );
  ND2S U18059 ( .I1(cnt_bdyn[2]), .I2(n30303), .O(n21153) );
  ND2S U18060 ( .I1(n30424), .I2(n30330), .O(n21151) );
  ND2S U18061 ( .I1(cnt_bdyn[3]), .I2(n30299), .O(n21145) );
  ND2S U18062 ( .I1(cnt_bdyn[2]), .I2(n30135), .O(n21147) );
  ND2S U18063 ( .I1(n30135), .I2(n30365), .O(n21146) );
  ND2S U18064 ( .I1(n30298), .I2(n30330), .O(n21114) );
  ND2S U18065 ( .I1(n30298), .I2(n30322), .O(n22811) );
  ND2 U18066 ( .I1(n16052), .I2(n18478), .O(n18884) );
  MAO222S U18067 ( .A1(gray_img[132]), .B1(n23438), .C1(n23437), .O(n23439) );
  MAO222S U18068 ( .A1(gray_img[131]), .B1(n23436), .C1(n23435), .O(n23437) );
  MAO222S U18069 ( .A1(gray_img[130]), .B1(n23434), .C1(n23433), .O(n23435) );
  AO22S U18070 ( .A1(n23462), .A2(n23458), .B1(n23446), .B2(n15982), .O(n15970) );
  OR2S U18071 ( .I1(n23462), .I2(n23458), .O(n15982) );
  MAO222 U18072 ( .A1(n23463), .B1(n23467), .C1(n23445), .O(n23446) );
  MAO222S U18073 ( .A1(n30119), .B1(n23482), .C1(n23478), .O(n23445) );
  ND2 U18074 ( .I1(n30383), .I2(n16010), .O(n18455) );
  ND2S U18075 ( .I1(n24407), .I2(n24400), .O(n24484) );
  OR2S U18076 ( .I1(n24795), .I2(n24794), .O(n24835) );
  AOI12HS U18077 ( .B1(n24331), .B2(n24294), .A1(n24293), .O(n24439) );
  ND3 U18078 ( .I1(n24464), .I2(n24463), .I3(n24462), .O(n24828) );
  AO12S U18079 ( .B1(n24382), .B2(n24647), .A1(n24360), .O(n24453) );
  INV1S U18080 ( .I(n24359), .O(n24454) );
  AO12S U18081 ( .B1(n24382), .B2(n24689), .A1(n24371), .O(n24495) );
  OR2S U18082 ( .I1(n24687), .I2(n24693), .O(n24692) );
  OR2S U18083 ( .I1(n24688), .I2(n24695), .O(n24691) );
  OA112 U18084 ( .C1(n24620), .C2(n24587), .A1(n24586), .B1(n24585), .O(n24790) );
  AO12S U18085 ( .B1(n24382), .B2(n24697), .A1(n24381), .O(n24508) );
  AOI12HS U18086 ( .B1(n24331), .B2(n24319), .A1(n24318), .O(n24507) );
  OR2S U18087 ( .I1(n24694), .I2(n24693), .O(n24701) );
  OR2S U18088 ( .I1(n24696), .I2(n24695), .O(n24700) );
  OA112 U18089 ( .C1(n24620), .C2(n24596), .A1(n24595), .B1(n24594), .O(n24785) );
  ND2S U18090 ( .I1(n24855), .I2(n24796), .O(n24800) );
  ND2S U18091 ( .I1(n24942), .I2(n19397), .O(n19403) );
  ND2 U18092 ( .I1(medfilt_state[2]), .I2(medfilt_state[1]), .O(n19087) );
  OR2S U18093 ( .I1(n30445), .I2(n30447), .O(n15975) );
  OA12S U18094 ( .B1(gray_scale_1[4]), .B2(n19944), .A1(n19943), .O(n19949) );
  ND2S U18095 ( .I1(gray_scale_1[3]), .I2(n30442), .O(n19947) );
  ND2S U18096 ( .I1(n18453), .I2(n18152), .O(n30359) );
  OAI12HS U18097 ( .B1(n17575), .B2(n17574), .A1(n17573), .O(n17577) );
  ND2S U18098 ( .I1(n17942), .I2(n17940), .O(n17573) );
  XNR2HS U18099 ( .I1(n17942), .I2(n17941), .O(n17946) );
  FA1S U18100 ( .A(n17897), .B(n17896), .CI(n17895), .CO(n17914), .S(n17907)
         );
  HA1S U18101 ( .A(cro_mac[2]), .B(n17881), .C(n17879), .S(n17888) );
  HA1S U18102 ( .A(cro_mac[1]), .B(n17885), .C(n17882), .S(n17887) );
  ND3S U18103 ( .I1(n16113), .I2(n25045), .I3(n25037), .O(n16086) );
  ND2S U18104 ( .I1(n25040), .I2(n24897), .O(n17950) );
  MAO222S U18105 ( .A1(n26552), .B1(gray_img[1556]), .C1(n26551), .O(n26553)
         );
  OR2S U18106 ( .I1(n24083), .I2(n24119), .O(n24086) );
  AN3S U18107 ( .I1(n24664), .I2(n24663), .I3(n24662), .O(n15984) );
  OR2S U18108 ( .I1(n24659), .I2(n24693), .O(n24664) );
  OR2S U18109 ( .I1(n24660), .I2(n24695), .O(n24663) );
  OR2S U18110 ( .I1(n21159), .I2(n21158), .O(n22487) );
  ND2S U18111 ( .I1(n21125), .I2(n30298), .O(n22853) );
  INV1S U18112 ( .I(n21933), .O(n22695) );
  INV1S U18113 ( .I(n22156), .O(n22810) );
  NR2 U18114 ( .I1(n18822), .I2(n18821), .O(n25282) );
  NR2 U18115 ( .I1(n18821), .I2(n25052), .O(n25244) );
  NR2 U18116 ( .I1(n18884), .I2(n25052), .O(n25193) );
  NR2 U18117 ( .I1(n18821), .I2(n24973), .O(n25085) );
  NR2 U18118 ( .I1(n18884), .I2(n24973), .O(n25272) );
  NR2 U18119 ( .I1(n24999), .I2(n18821), .O(n25325) );
  NR2 U18120 ( .I1(n18822), .I2(n24998), .O(n19406) );
  NR2 U18121 ( .I1(n25052), .I2(n24998), .O(n19844) );
  NR2 U18122 ( .I1(n24973), .I2(n24998), .O(n25351) );
  NR2 U18123 ( .I1(n24973), .I2(n25051), .O(n25355) );
  NR2 U18124 ( .I1(n24999), .I2(n24998), .O(n25365) );
  AN2S U18125 ( .I1(n18383), .I2(n24903), .O(n18392) );
  OR2S U18126 ( .I1(n21114), .I2(n21146), .O(n22865) );
  NR2 U18127 ( .I1(n18884), .I2(n24999), .O(n25216) );
  OA12S U18128 ( .B1(cnt[0]), .B2(n18403), .A1(n18418), .O(n30400) );
  ND3S U18129 ( .I1(n30321), .I2(n30353), .I3(n30323), .O(n30129) );
  INV1S U18130 ( .I(n18455), .O(n18642) );
  OR2S U18131 ( .I1(n16089), .I2(cs[2]), .O(n24910) );
  ND2S U18132 ( .I1(n30303), .I2(n30365), .O(n30306) );
  OR2S U18133 ( .I1(n24485), .I2(n24484), .O(n24894) );
  OR2S U18134 ( .I1(cnt_cro_3[1]), .I2(cnt_cro_3[0]), .O(n24939) );
  INV1S U18135 ( .I(n24819), .O(n24885) );
  ND3 U18136 ( .I1(n24483), .I2(n24482), .I3(n24481), .O(n24887) );
  BUF2 U18137 ( .I(n19087), .O(n24919) );
  OR2S U18138 ( .I1(image_size_reg_set[1]), .I2(image_size_reg_set[0]), .O(
        n24901) );
  AN2S U18139 ( .I1(cnt_bdyn[5]), .I2(n30356), .O(n30358) );
  FA1S U18140 ( .A(image[1]), .B(gray_scale_1[1]), .CI(n30347), .CO(n30345), 
        .S(n30348) );
  FA1S U18141 ( .A(image[2]), .B(gray_scale_1[2]), .CI(n30345), .CO(n30343), 
        .S(n30346) );
  FA1S U18142 ( .A(image[3]), .B(gray_scale_1[3]), .CI(n30343), .CO(n30341), 
        .S(n30344) );
  ND2S U18143 ( .I1(n30349), .I2(gray_scale_0[7]), .O(n23055) );
  MAO222 U18144 ( .A1(n30338), .B1(gray_scale_0[6]), .C1(n23053), .O(n23054)
         );
  MAO222 U18145 ( .A1(n30421), .B1(gray_scale_0[5]), .C1(n23052), .O(n23053)
         );
  INV1S U18146 ( .I(image[1]), .O(n30415) );
  OA12 U18147 ( .B1(gray_scale_0[7]), .B2(n30423), .A1(n30422), .O(n30419) );
  ND2S U18148 ( .I1(cnt_dyn[0]), .I2(cnt_dyn[1]), .O(n30251) );
  OR2S U18149 ( .I1(cnt_cro_3[1]), .I2(n16090), .O(n24943) );
  ND2S U18150 ( .I1(n24942), .I2(n25040), .O(n24944) );
  OR2S U18151 ( .I1(cs[1]), .I2(n24910), .O(n30390) );
  ND2S U18152 ( .I1(n17993), .I2(cro_mac[15]), .O(n18038) );
  ND2S U18153 ( .I1(n17992), .I2(n17991), .O(n18047) );
  OR2S U18154 ( .I1(n17888), .I2(n17889), .O(n30206) );
  ND2S U18155 ( .I1(n30135), .I2(n30133), .O(n30143) );
  ND2S U18156 ( .I1(n30134), .I2(n30135), .O(n30144) );
  ND2S U18157 ( .I1(n30136), .I2(n30135), .O(n30145) );
  ND2S U18158 ( .I1(n30303), .I2(n30133), .O(n30138) );
  ND2S U18159 ( .I1(n30134), .I2(n30303), .O(n30137) );
  ND2S U18160 ( .I1(n30136), .I2(n30303), .O(n30139) );
  MUX2S U18161 ( .A(n30056), .B(n28581), .S(gray_img[672]), .O(n23539) );
  MUX2S U18162 ( .A(gray_img[473]), .B(gray_img[345]), .S(n27353), .O(n26823)
         );
  MUX2S U18163 ( .A(gray_img[1972]), .B(gray_img[1844]), .S(n23162), .O(n23178) );
  MUX2S U18164 ( .A(gray_img[1628]), .B(gray_img[1756]), .S(n25577), .O(n25559) );
  MUX2S U18165 ( .A(gray_img[1684]), .B(gray_img[1556]), .S(n29577), .O(n29536) );
  MUX2S U18166 ( .A(gray_img[1156]), .B(gray_img[1028]), .S(n29731), .O(n29716) );
  MUX2S U18167 ( .A(gray_img[212]), .B(gray_img[84]), .S(n23483), .O(n16046)
         );
  ND2S U18168 ( .I1(n28530), .I2(n26842), .O(n16058) );
  MUX2S U18169 ( .A(gray_img[1685]), .B(gray_img[1557]), .S(n29577), .O(n29531) );
  MUX2S U18170 ( .A(gray_img[477]), .B(gray_img[349]), .S(n27353), .O(n26803)
         );
  MUX2S U18171 ( .A(gray_img[1973]), .B(gray_img[1845]), .S(n23162), .O(n23183) );
  MUX2S U18172 ( .A(gray_img[1974]), .B(gray_img[1846]), .S(n23162), .O(n23188) );
  MUX2S U18173 ( .A(gray_img[1630]), .B(gray_img[1758]), .S(n25577), .O(n25549) );
  MUX2S U18174 ( .A(gray_img[1486]), .B(gray_img[1358]), .S(n23536), .O(n23544) );
  INV1 U18175 ( .I(n16006), .O(n29427) );
  AN2S U18176 ( .I1(n19127), .I2(medfilt_out_reg[6]), .O(n18097) );
  ND2S U18177 ( .I1(n30132), .I2(n30133), .O(n30141) );
  ND2S U18178 ( .I1(n30134), .I2(n30132), .O(n30140) );
  ND2S U18179 ( .I1(n30136), .I2(n30132), .O(n30142) );
  ND2S U18180 ( .I1(n30329), .I2(n30301), .O(n30335) );
  AO12S U18181 ( .B1(n30012), .B2(n29970), .A1(n29969), .O(n13735) );
  ND2S U18182 ( .I1(n15885), .I2(n30006), .O(n29966) );
  MUX2S U18183 ( .A(n30005), .B(n30006), .S(gray_img[257]), .O(n29967) );
  AO12S U18184 ( .B1(n29604), .B2(n29592), .A1(n29591), .O(n13686) );
  ND2S U18185 ( .I1(n15933), .I2(n29598), .O(n29588) );
  MUX2S U18186 ( .A(n29587), .B(n29598), .S(gray_img[905]), .O(n29589) );
  ND2S U18187 ( .I1(n28806), .I2(n23241), .O(n23245) );
  MUX2S U18188 ( .A(n29587), .B(n28807), .S(gray_img[401]), .O(n23243) );
  AO12S U18189 ( .B1(n15886), .B2(n27261), .A1(n27191), .O(n14411) );
  MUX2S U18190 ( .A(n28534), .B(n27259), .S(gray_img[969]), .O(n27191) );
  ND2S U18191 ( .I1(n19755), .I2(n19754), .O(n14260) );
  MUX2S U18192 ( .A(n27447), .B(n26757), .S(gray_img[344]), .O(n26752) );
  ND2S U18193 ( .I1(n15884), .I2(n20389), .O(n18902) );
  MUX2S U18194 ( .A(n29566), .B(n20389), .S(gray_img[1937]), .O(n18903) );
  ND2S U18195 ( .I1(n15884), .I2(n20843), .O(n20844) );
  MUX2S U18196 ( .A(n20842), .B(n20843), .S(gray_img[1313]), .O(n20845) );
  ND2S U18197 ( .I1(n15884), .I2(n20379), .O(n18507) );
  MUX2S U18198 ( .A(n29587), .B(n20379), .S(gray_img[1185]), .O(n18508) );
  MUX2S U18199 ( .A(n20842), .B(n20509), .S(gray_img[1656]), .O(n19175) );
  AO12S U18200 ( .B1(n15886), .B2(n26224), .A1(n26223), .O(n14416) );
  AO12S U18201 ( .B1(n26939), .B2(n26938), .A1(n26937), .O(n14212) );
  ND2S U18202 ( .I1(n15885), .I2(n26932), .O(n26933) );
  MUX2S U18203 ( .A(n29032), .B(n26932), .S(gray_img[161]), .O(n26934) );
  MUX2S U18204 ( .A(n29597), .B(n20881), .S(gray_img[1537]), .O(n20878) );
  AO12S U18205 ( .B1(n27121), .B2(n27113), .A1(n27112), .O(n13781) );
  MUX2S U18206 ( .A(n29566), .B(n27114), .S(gray_img[296]), .O(n27110) );
  AO12S U18207 ( .B1(n27121), .B2(n27120), .A1(n27119), .O(n14159) );
  ND2S U18208 ( .I1(n15885), .I2(n27114), .O(n27115) );
  MUX2S U18209 ( .A(n30044), .B(n27114), .S(gray_img[297]), .O(n27116) );
  AO12S U18210 ( .B1(n27556), .B2(n27542), .A1(n27541), .O(n14238) );
  ND2S U18211 ( .I1(n15933), .I2(n27550), .O(n27538) );
  MUX2S U18212 ( .A(n29032), .B(n27550), .S(gray_img[49]), .O(n27539) );
  AO12S U18213 ( .B1(n30012), .B2(n30011), .A1(n30010), .O(n13736) );
  ND3S U18214 ( .I1(n30009), .I2(n30008), .I3(n30007), .O(n30010) );
  AO12S U18215 ( .B1(n28214), .B2(n28133), .A1(n28132), .O(n13697) );
  ND2S U18216 ( .I1(n15928), .I2(n28208), .O(n28129) );
  MUX2S U18217 ( .A(n30005), .B(n28208), .S(gray_img[689]), .O(n28130) );
  AO12S U18218 ( .B1(n30038), .B2(n29386), .A1(n29385), .O(n14271) );
  ND2S U18219 ( .I1(n15931), .I2(n30032), .O(n29382) );
  MUX2S U18220 ( .A(n30050), .B(n30032), .S(gray_img[393]), .O(n29383) );
  AO12S U18221 ( .B1(n29040), .B2(n29016), .A1(n29015), .O(n13728) );
  AO12S U18222 ( .B1(n28459), .B2(n28431), .A1(n28430), .O(n13741) );
  AO12S U18223 ( .B1(n29040), .B2(n29039), .A1(n29038), .O(n13966) );
  ND2S U18224 ( .I1(n15885), .I2(n29033), .O(n29034) );
  MUX2S U18225 ( .A(n29032), .B(n29033), .S(gray_img[657]), .O(n29035) );
  AO12S U18226 ( .B1(n30109), .B2(n30017), .A1(n30016), .O(n14272) );
  ND2S U18227 ( .I1(n15933), .I2(n30103), .O(n30013) );
  MUX2S U18228 ( .A(n15904), .B(n30103), .S(gray_img[385]), .O(n30014) );
  AO12S U18229 ( .B1(n26473), .B2(n26444), .A1(n26443), .O(n13763) );
  MUX2S U18230 ( .A(n30056), .B(n26466), .S(gray_img[440]), .O(n26441) );
  AO12S U18231 ( .B1(n28459), .B2(n28458), .A1(n28457), .O(n14027) );
  ND2S U18232 ( .I1(n15885), .I2(n28452), .O(n28453) );
  MUX2S U18233 ( .A(n29032), .B(n28452), .S(gray_img[553]), .O(n28454) );
  AO12S U18234 ( .B1(n25619), .B2(n25618), .A1(n25617), .O(n13682) );
  ND2S U18235 ( .I1(n15931), .I2(n25612), .O(n25613) );
  MUX2S U18236 ( .A(n30044), .B(n25612), .S(gray_img[937]), .O(n25614) );
  AO12S U18237 ( .B1(n26473), .B2(n26472), .A1(n26471), .O(n14097) );
  ND2S U18238 ( .I1(n15933), .I2(n26466), .O(n26467) );
  MUX2S U18239 ( .A(n15904), .B(n26466), .S(gray_img[441]), .O(n26468) );
  OA12S U18240 ( .B1(n29884), .B2(n28709), .A1(n28708), .O(n28710) );
  MUX2S U18241 ( .A(n15904), .B(n28707), .S(gray_img[273]), .O(n28708) );
  AO12S U18242 ( .B1(n27692), .B2(n27664), .A1(n27663), .O(n13793) );
  MUX2S U18243 ( .A(n30050), .B(n27685), .S(gray_img[184]), .O(n27661) );
  AO12S U18244 ( .B1(n26489), .B2(n26478), .A1(n26477), .O(n14141) );
  ND2S U18245 ( .I1(n15933), .I2(n26483), .O(n26474) );
  MUX2S U18246 ( .A(n15904), .B(n26483), .S(gray_img[313]), .O(n26475) );
  AO12S U18247 ( .B1(n27692), .B2(n27691), .A1(n27690), .O(n14185) );
  ND2S U18248 ( .I1(n15885), .I2(n27685), .O(n27686) );
  MUX2S U18249 ( .A(n30050), .B(n27685), .S(gray_img[185]), .O(n27687) );
  AO12S U18250 ( .B1(n30098), .B2(n29492), .A1(n29491), .O(n13687) );
  ND2S U18251 ( .I1(n15933), .I2(n30092), .O(n29488) );
  MUX2S U18252 ( .A(n29597), .B(n30092), .S(gray_img[897]), .O(n29489) );
  AO12S U18253 ( .B1(n26849), .B2(n26848), .A1(n26847), .O(n14247) );
  MUX2S U18254 ( .A(n30044), .B(n26842), .S(gray_img[41]), .O(n26844) );
  AO12S U18255 ( .B1(n27378), .B2(n27370), .A1(n27369), .O(n13802) );
  AO12S U18256 ( .B1(n27378), .B2(n27377), .A1(n27376), .O(n13801) );
  ND2S U18257 ( .I1(n15885), .I2(n27371), .O(n27372) );
  MUX2S U18258 ( .A(n30050), .B(n27371), .S(gray_img[17]), .O(n27373) );
  ND2S U18259 ( .I1(n30120), .I2(n23478), .O(n23481) );
  AO12S U18260 ( .B1(n28128), .B2(n28127), .A1(n28126), .O(n14018) );
  ND2S U18261 ( .I1(n15933), .I2(n28121), .O(n28122) );
  MUX2S U18262 ( .A(n29597), .B(n28121), .S(gray_img[561]), .O(n28123) );
  ND2S U18263 ( .I1(n30020), .I2(n29193), .O(n29196) );
  OA12S U18264 ( .B1(n29884), .B2(n30023), .A1(n29194), .O(n29195) );
  MUX2S U18265 ( .A(n30056), .B(n30021), .S(gray_img[913]), .O(n29194) );
  AO12S U18266 ( .B1(n28588), .B2(n28587), .A1(n28586), .O(n13699) );
  ND2S U18267 ( .I1(n15933), .I2(n28581), .O(n28582) );
  MUX2S U18268 ( .A(n30044), .B(n28581), .S(gray_img[673]), .O(n28583) );
  ND2S U18269 ( .I1(n23492), .I2(n23367), .O(n23370) );
  MUX2S U18270 ( .A(n30050), .B(n23493), .S(gray_img[569]), .O(n23368) );
  ND2S U18271 ( .I1(n23492), .I2(n23491), .O(n23497) );
  MUX2S U18272 ( .A(n30044), .B(n23493), .S(gray_img[568]), .O(n23494) );
  ND2S U18273 ( .I1(n29993), .I2(n29706), .O(n29709) );
  OA12S U18274 ( .B1(n29884), .B2(n29996), .A1(n29707), .O(n29708) );
  MUX2S U18275 ( .A(n15904), .B(n29994), .S(gray_img[641]), .O(n29707) );
  ND2S U18276 ( .I1(n28727), .I2(n28241), .O(n28244) );
  OA12S U18277 ( .B1(n29884), .B2(n28730), .A1(n28242), .O(n28243) );
  MUX2S U18278 ( .A(n15904), .B(n28728), .S(gray_img[409]), .O(n28242) );
  ND2S U18279 ( .I1(n23121), .I2(n23120), .O(n23125) );
  MUX2S U18280 ( .A(n29566), .B(n25151), .S(gray_img[425]), .O(n23122) );
  ND2S U18281 ( .I1(n26327), .I2(n26318), .O(n26319) );
  OA12S U18282 ( .B1(n29884), .B2(n26324), .A1(n26317), .O(n26320) );
  MUX2S U18283 ( .A(n15904), .B(n26322), .S(gray_img[305]), .O(n26317) );
  ND2S U18284 ( .I1(n26327), .I2(n26326), .O(n26328) );
  OA12S U18285 ( .B1(n29734), .B2(n26324), .A1(n26323), .O(n26329) );
  OA12S U18286 ( .B1(n29734), .B2(n25607), .A1(n25579), .O(n25580) );
  OA12S U18287 ( .B1(n29884), .B2(n29742), .A1(n29741), .O(n29743) );
  MUX2S U18288 ( .A(n15904), .B(n29740), .S(gray_img[513]), .O(n29741) );
  OA12S U18289 ( .B1(n29734), .B2(n29742), .A1(n29733), .O(n29735) );
  ND2S U18290 ( .I1(n29043), .I2(n23044), .O(n23047) );
  MUX2S U18291 ( .A(n30050), .B(n29044), .S(gray_img[530]), .O(n23045) );
  ND2S U18292 ( .I1(n19781), .I2(n19780), .O(n14088) );
  MUX2S U18293 ( .A(n29566), .B(n20255), .S(gray_img[1040]), .O(n19780) );
  MUX2S U18294 ( .A(n30044), .B(n20392), .S(gray_img[1280]), .O(n19318) );
  MUX2S U18295 ( .A(n29566), .B(n20836), .S(gray_img[1320]), .O(n19346) );
  MUX2S U18296 ( .A(n29587), .B(n20296), .S(gray_img[1816]), .O(n19338) );
  ND2S U18297 ( .I1(n15884), .I2(n20354), .O(n20355) );
  MUX2S U18298 ( .A(n29597), .B(n20354), .S(gray_img[1809]), .O(n20356) );
  AO12S U18299 ( .B1(n15886), .B2(n26942), .A1(n26862), .O(n14443) );
  MUX2S U18300 ( .A(n28534), .B(n26940), .S(gray_img[457]), .O(n26862) );
  AO12S U18301 ( .B1(n15886), .B2(n27829), .A1(n26225), .O(n14408) );
  AO12S U18302 ( .B1(n15886), .B2(n28560), .A1(n28537), .O(n14347) );
  MUX2S U18303 ( .A(n27447), .B(n28558), .S(gray_img[1481]), .O(n28537) );
  AO12S U18304 ( .B1(n15886), .B2(n26726), .A1(n26710), .O(n14457) );
  AO12S U18305 ( .B1(n15886), .B2(n27013), .A1(n27010), .O(n14434) );
  MUX2S U18306 ( .A(n28534), .B(n27011), .S(gray_img[593]), .O(n27010) );
  MUX2S U18307 ( .A(n30056), .B(n20362), .S(gray_img[1296]), .O(n19108) );
  MUX2S U18308 ( .A(n29597), .B(n20862), .S(gray_img[1840]), .O(n19114) );
  ND2S U18309 ( .I1(n20636), .I2(n20635), .O(n14420) );
  ND2S U18310 ( .I1(n15884), .I2(n20634), .O(n20636) );
  ND2S U18311 ( .I1(n19837), .I2(n19836), .O(n14431) );
  MUX2S U18312 ( .A(n20274), .B(n20830), .S(intadd_103_CI), .O(n19836) );
  ND2S U18313 ( .I1(n20633), .I2(n20632), .O(n14460) );
  ND2S U18314 ( .I1(n15886), .I2(n20631), .O(n20633) );
  MUX2S U18315 ( .A(n30044), .B(n20631), .S(gray_img[193]), .O(n20632) );
  ND2S U18316 ( .I1(n19925), .I2(n19924), .O(n14266) );
  ND2S U18317 ( .I1(n19906), .I2(n19905), .O(n14468) );
  ND2S U18318 ( .I1(n20625), .I2(n20624), .O(n14428) );
  ND2S U18319 ( .I1(n15928), .I2(n20623), .O(n20625) );
  MUX2S U18320 ( .A(n29587), .B(n20623), .S(gray_img[705]), .O(n20624) );
  ND2S U18321 ( .I1(n19785), .I2(n19784), .O(n14402) );
  ND2S U18322 ( .I1(n15886), .I2(n20255), .O(n19785) );
  MUX2S U18323 ( .A(n29597), .B(n20255), .S(gray_img[1041]), .O(n19784) );
  ND2S U18324 ( .I1(n19884), .I2(n19883), .O(n14444) );
  ND2S U18325 ( .I1(n15884), .I2(n20483), .O(n19884) );
  ND2S U18326 ( .I1(n19890), .I2(n19889), .O(n14645) );
  ND2S U18327 ( .I1(n15883), .I2(n20483), .O(n19890) );
  ND2S U18328 ( .I1(n19730), .I2(n19729), .O(n14462) );
  MUX2S U18329 ( .A(n30050), .B(n20499), .S(gray_img[113]), .O(n19729) );
  ND2S U18330 ( .I1(n19716), .I2(n19715), .O(n14454) );
  MUX2S U18331 ( .A(n30056), .B(n20260), .S(gray_img[241]), .O(n19715) );
  ND2S U18332 ( .I1(n19745), .I2(n19744), .O(n14083) );
  MUX2S U18333 ( .A(n30056), .B(n20760), .S(gray_img[1080]), .O(n19744) );
  MUX2S U18334 ( .A(n27447), .B(n26877), .S(gray_img[72]), .O(n26872) );
  AO12S U18335 ( .B1(n19092), .B2(n26722), .A1(n26715), .O(n14264) );
  MUX2S U18336 ( .A(n28534), .B(n26720), .S(gray_img[80]), .O(n26715) );
  ND2S U18337 ( .I1(n15884), .I2(n20608), .O(n20610) );
  ND2S U18338 ( .I1(n15932), .I2(n20614), .O(n20616) );
  ND2S U18339 ( .I1(n15884), .I2(n20591), .O(n20592) );
  MUX2S U18340 ( .A(n29587), .B(n20591), .S(gray_img[577]), .O(n20593) );
  ND2S U18341 ( .I1(n15885), .I2(n20565), .O(n20567) );
  MUX2S U18342 ( .A(n30005), .B(n20565), .S(gray_img[633]), .O(n20566) );
  ND2S U18343 ( .I1(n15933), .I2(n20528), .O(n20530) );
  ND2S U18344 ( .I1(n15885), .I2(n20504), .O(n20506) );
  MUX2S U18345 ( .A(n30056), .B(n20504), .S(gray_img[1857]), .O(n20505) );
  AO12S U18346 ( .B1(n15884), .B2(n26722), .A1(n26721), .O(n14466) );
  MUX2S U18347 ( .A(n28534), .B(n26720), .S(gray_img[81]), .O(n26721) );
  AO12S U18348 ( .B1(n15886), .B2(n26747), .A1(n26740), .O(n14442) );
  AO12S U18349 ( .B1(n15886), .B2(n25778), .A1(n25777), .O(n14312) );
  MUX2S U18350 ( .A(n15889), .B(n26741), .S(gray_img[336]), .O(n26742) );
  MUX2S U18351 ( .A(n27447), .B(n25830), .S(gray_img[1888]), .O(n25831) );
  AO12S U18352 ( .B1(n15886), .B2(n27009), .A1(n27008), .O(n14426) );
  MUX2S U18353 ( .A(n27447), .B(n27007), .S(gray_img[721]), .O(n27008) );
  AO12S U18354 ( .B1(n15886), .B2(n28596), .A1(n28343), .O(n14362) );
  MUX2S U18355 ( .A(n27447), .B(n28594), .S(gray_img[1361]), .O(n28343) );
  AO12S U18356 ( .B1(n15886), .B2(n28342), .A1(n28341), .O(n14346) );
  MUX2S U18357 ( .A(n27447), .B(n28340), .S(gray_img[1489]), .O(n28341) );
  AO12S U18358 ( .B1(n15886), .B2(n26709), .A1(n26708), .O(n14465) );
  MUX2S U18359 ( .A(n27447), .B(n26707), .S(gray_img[89]), .O(n26708) );
  AO12S U18360 ( .B1(n15886), .B2(n27243), .A1(n27134), .O(n14427) );
  AO12S U18361 ( .B1(n15886), .B2(n26996), .A1(n26995), .O(n14425) );
  MUX2S U18362 ( .A(n29587), .B(n20605), .S(gray_img[1681]), .O(n19617) );
  ND2S U18363 ( .I1(n15884), .I2(n20746), .O(n20673) );
  MUX2S U18364 ( .A(n29566), .B(n20746), .S(gray_img[1977]), .O(n20672) );
  ND2S U18365 ( .I1(n15937), .I2(n20746), .O(n20715) );
  MUX2S U18366 ( .A(n29566), .B(n20746), .S(gray_img[1978]), .O(n20714) );
  ND2S U18367 ( .I1(n15932), .I2(n20740), .O(n20701) );
  MUX2S U18368 ( .A(n29597), .B(n20740), .S(gray_img[1849]), .O(n20700) );
  ND2S U18369 ( .I1(n15884), .I2(n20695), .O(n20681) );
  MUX2S U18370 ( .A(n30056), .B(n20695), .S(gray_img[1337]), .O(n20680) );
  ND2S U18371 ( .I1(n27512), .I2(n20737), .O(n20638) );
  MUX2S U18372 ( .A(n30044), .B(n20737), .S(gray_img[1721]), .O(n20637) );
  ND2S U18373 ( .I1(n27512), .I2(n20709), .O(n20677) );
  MUX2S U18374 ( .A(n20830), .B(n20709), .S(gray_img[1465]), .O(n20676) );
  ND2S U18375 ( .I1(n15928), .I2(n20836), .O(n20837) );
  MUX2S U18376 ( .A(n29566), .B(n20836), .S(gray_img[1321]), .O(n20838) );
  ND2S U18377 ( .I1(n15885), .I2(n20814), .O(n20775) );
  MUX2S U18378 ( .A(n29566), .B(n20814), .S(gray_img[1449]), .O(n20776) );
  ND2S U18379 ( .I1(n27512), .I2(n20827), .O(n20769) );
  MUX2S U18380 ( .A(n30050), .B(n20827), .S(gray_img[1705]), .O(n20770) );
  MUX2S U18381 ( .A(n29566), .B(n20583), .S(gray_img[1665]), .O(n19557) );
  ND2S U18382 ( .I1(n15930), .I2(n20373), .O(n18881) );
  MUX2S U18383 ( .A(n20842), .B(n20373), .S(gray_img[1921]), .O(n18882) );
  ND2S U18384 ( .I1(n27512), .I2(n20392), .O(n18874) );
  MUX2S U18385 ( .A(n30050), .B(n20392), .S(gray_img[1281]), .O(n18875) );
  ND2S U18386 ( .I1(n27512), .I2(n20359), .O(n18866) );
  ND2S U18387 ( .I1(n15930), .I2(n20811), .O(n20809) );
  MUX2S U18388 ( .A(n20808), .B(n20811), .S(gray_img[1441]), .O(n20810) );
  ND2S U18389 ( .I1(n15928), .I2(n20846), .O(n20767) );
  MUX2S U18390 ( .A(n30050), .B(n20846), .S(gray_img[1713]), .O(n20768) );
  ND2S U18391 ( .I1(n15932), .I2(n20862), .O(n20763) );
  MUX2S U18392 ( .A(n29597), .B(n20862), .S(gray_img[1841]), .O(n20764) );
  ND2S U18393 ( .I1(n15884), .I2(n20849), .O(n20765) );
  MUX2S U18394 ( .A(n29597), .B(n20849), .S(gray_img[1969]), .O(n20766) );
  ND2S U18395 ( .I1(n15884), .I2(n20787), .O(n20788) );
  MUX2S U18396 ( .A(n30056), .B(n20787), .S(gray_img[1697]), .O(n20789) );
  ND2S U18397 ( .I1(n15885), .I2(n20743), .O(n20708) );
  MUX2S U18398 ( .A(n29587), .B(n20743), .S(gray_img[1089]), .O(n20707) );
  ND2S U18399 ( .I1(n15884), .I2(n20716), .O(n20679) );
  MUX2S U18400 ( .A(n30050), .B(n20716), .S(gray_img[1145]), .O(n20678) );
  ND2S U18401 ( .I1(n15885), .I2(n20702), .O(n20704) );
  MUX2S U18402 ( .A(n30056), .B(n20702), .S(gray_img[1217]), .O(n20703) );
  ND2S U18403 ( .I1(n15932), .I2(n20655), .O(n20657) );
  MUX2S U18404 ( .A(n20808), .B(n20655), .S(gray_img[1273]), .O(n20656) );
  ND2S U18405 ( .I1(n15885), .I2(n20728), .O(n20688) );
  MUX2S U18406 ( .A(n20808), .B(n20728), .S(gray_img[1129]), .O(n20687) );
  ND2S U18407 ( .I1(n15931), .I2(n20719), .O(n20721) );
  MUX2S U18408 ( .A(n20842), .B(n20719), .S(gray_img[1257]), .O(n20720) );
  MUX2S U18409 ( .A(n29587), .B(n20553), .S(gray_img[1161]), .O(n19504) );
  ND2S U18410 ( .I1(n15884), .I2(n20427), .O(n18728) );
  MUX2S U18411 ( .A(n20842), .B(n20427), .S(gray_img[1289]), .O(n18727) );
  MUX2S U18412 ( .A(n30050), .B(n20553), .S(gray_img[1160]), .O(n19046) );
  ND2S U18413 ( .I1(n15884), .I2(n20440), .O(n19643) );
  MUX2S U18414 ( .A(n30050), .B(n20440), .S(gray_img[1513]), .O(n19642) );
  ND2S U18415 ( .I1(n15884), .I2(n20159), .O(n18639) );
  MUX2S U18416 ( .A(n29597), .B(n20159), .S(gray_img[1177]), .O(n18640) );
  ND2S U18417 ( .I1(n15883), .I2(n20159), .O(n18637) );
  MUX2S U18418 ( .A(n29597), .B(n20159), .S(gray_img[1178]), .O(n18638) );
  MUX2S U18419 ( .A(n29597), .B(n20184), .S(gray_img[1049]), .O(n19611) );
  MUX2S U18420 ( .A(n29587), .B(n20296), .S(gray_img[1817]), .O(n19619) );
  ND2S U18421 ( .I1(n15884), .I2(n19970), .O(n18801) );
  MUX2S U18422 ( .A(n30005), .B(n19970), .S(gray_img[1945]), .O(n18802) );
  MUX2S U18423 ( .A(n20808), .B(n20719), .S(gray_img[1256]), .O(n19048) );
  MUX2S U18424 ( .A(n30005), .B(n20534), .S(gray_img[625]), .O(n19532) );
  MUX2S U18425 ( .A(n30005), .B(n20054), .S(gray_img[753]), .O(n19530) );
  MUX2S U18426 ( .A(n15904), .B(n20099), .S(gray_img[1017]), .O(n19518) );
  ND2S U18427 ( .I1(n15884), .I2(n20209), .O(n18947) );
  MUX2S U18428 ( .A(n29587), .B(n20684), .S(gray_img[1472]), .O(n19170) );
  MUX2S U18429 ( .A(n29587), .B(n20580), .S(gray_img[960]), .O(n19032) );
  AO12S U18430 ( .B1(n15886), .B2(n26879), .A1(n26878), .O(n14467) );
  MUX2S U18431 ( .A(n27447), .B(n26877), .S(gray_img[73]), .O(n26878) );
  AO12S U18432 ( .B1(n15886), .B2(n27545), .A1(n27391), .O(n14464) );
  MUX2S U18433 ( .A(n27447), .B(n27543), .S(gray_img[97]), .O(n27391) );
  AO12S U18434 ( .B1(n15886), .B2(n26759), .A1(n26758), .O(n14449) );
  MUX2S U18435 ( .A(n27447), .B(n26757), .S(gray_img[345]), .O(n26758) );
  AO12S U18436 ( .B1(n15886), .B2(n27352), .A1(n26760), .O(n14441) );
  MUX2S U18437 ( .A(n27447), .B(n27350), .S(gray_img[473]), .O(n26760) );
  MUX2S U18438 ( .A(n29587), .B(n20480), .S(gray_img[488]), .O(n19824) );
  ND2S U18439 ( .I1(n15884), .I2(n20235), .O(n19423) );
  MUX2S U18440 ( .A(n29597), .B(n20235), .S(gray_img[1033]), .O(n19422) );
  MUX2S U18441 ( .A(n29597), .B(n20235), .S(gray_img[1034]), .O(n19648) );
  MUX2S U18442 ( .A(n29587), .B(n20611), .S(gray_img[1064]), .O(n19676) );
  ND2S U18443 ( .I1(n15884), .I2(n20611), .O(n19687) );
  MUX2S U18444 ( .A(n29587), .B(n20611), .S(gray_img[1065]), .O(n19686) );
  ND2S U18445 ( .I1(n15884), .I2(n20240), .O(n19713) );
  MUX2S U18446 ( .A(n29587), .B(n20240), .S(gray_img[1153]), .O(n19712) );
  ND2S U18447 ( .I1(n15883), .I2(n20316), .O(n19769) );
  MUX2S U18448 ( .A(n29566), .B(n20316), .S(gray_img[1170]), .O(n19768) );
  ND2S U18449 ( .I1(n15884), .I2(n20435), .O(n19681) );
  MUX2S U18450 ( .A(n29566), .B(n20435), .S(gray_img[1193]), .O(n19680) );
  ND2S U18451 ( .I1(n15884), .I2(n20124), .O(n19635) );
  MUX2S U18452 ( .A(n20808), .B(n20124), .S(gray_img[1137]), .O(n19634) );
  MUX2S U18453 ( .A(n29587), .B(n20063), .S(gray_img[1904]), .O(n19068) );
  ND2S U18454 ( .I1(n15884), .I2(n25942), .O(n18585) );
  ND2S U18455 ( .I1(n15884), .I2(n20522), .O(n18499) );
  MUX2S U18456 ( .A(n30044), .B(n20522), .S(gray_img[369]), .O(n18498) );
  MUX2S U18457 ( .A(n30056), .B(n20477), .S(gray_img[497]), .O(n19526) );
  AO12S U18458 ( .B1(n15886), .B2(n25836), .A1(n25833), .O(n14280) );
  AO12S U18459 ( .B1(n15886), .B2(n27390), .A1(n27389), .O(n14456) );
  MUX2S U18460 ( .A(n27447), .B(n27388), .S(gray_img[225]), .O(n27389) );
  AO12S U18461 ( .B1(n15886), .B2(n27449), .A1(n27441), .O(n14448) );
  AO12S U18462 ( .B1(n15886), .B2(n27774), .A1(n27450), .O(n14440) );
  MUX2S U18463 ( .A(n27447), .B(n27772), .S(gray_img[481]), .O(n27450) );
  AO12S U18464 ( .B1(n15886), .B2(n27105), .A1(n26997), .O(n14433) );
  MUX2S U18465 ( .A(n27447), .B(n27103), .S(gray_img[601]), .O(n26997) );
  AO12S U18466 ( .B1(n15885), .B2(n27069), .A1(n27066), .O(n14418) );
  AO12S U18467 ( .B1(n15883), .B2(n27069), .A1(n27062), .O(n14619) );
  AO12S U18468 ( .B1(n15885), .B2(n30065), .A1(n27082), .O(n14417) );
  AO12S U18469 ( .B1(n15937), .B2(n30065), .A1(n27078), .O(n14618) );
  AO12S U18470 ( .B1(n15885), .B2(n27065), .A1(n27064), .O(n14410) );
  AO12S U18471 ( .B1(n15885), .B2(n27081), .A1(n27080), .O(n14409) );
  AO12S U18472 ( .B1(n15885), .B2(n28031), .A1(n28030), .O(n14376) );
  AO12S U18473 ( .B1(n15885), .B2(n25899), .A1(n25779), .O(n14328) );
  MUX2S U18474 ( .A(n30044), .B(n20082), .S(gray_img[121]), .O(n19462) );
  MUX2S U18475 ( .A(n29566), .B(n20496), .S(gray_img[249]), .O(n19486) );
  MUX2S U18476 ( .A(n30044), .B(n20556), .S(gray_img[1529]), .O(n19490) );
  ND2S U18477 ( .I1(n15884), .I2(n20547), .O(n18792) );
  MUX2S U18478 ( .A(n30056), .B(n20430), .S(gray_img[1912]), .O(n18743) );
  ND2S U18479 ( .I1(n15884), .I2(n20430), .O(n18786) );
  MUX2S U18480 ( .A(n29566), .B(n20430), .S(gray_img[1913]), .O(n18785) );
  MUX2S U18481 ( .A(n30044), .B(n20716), .S(gray_img[1144]), .O(n18779) );
  OA12S U18482 ( .B1(n29884), .B2(n29046), .A1(n23373), .O(n23374) );
  ND2S U18483 ( .I1(n29043), .I2(n23372), .O(n23375) );
  MUX2S U18484 ( .A(n30050), .B(n29044), .S(gray_img[529]), .O(n23373) );
  ND2S U18485 ( .I1(n15884), .I2(n20857), .O(n20858) );
  MUX2S U18486 ( .A(n30044), .B(n20857), .S(gray_img[1201]), .O(n20859) );
  ND2S U18487 ( .I1(n20750), .I2(n20749), .O(n14381) );
  ND2S U18488 ( .I1(n15884), .I2(n20757), .O(n20750) );
  MUX2S U18489 ( .A(n30044), .B(n20757), .S(gray_img[1209]), .O(n20749) );
  ND2S U18490 ( .I1(n15884), .I2(n20376), .O(n18876) );
  MUX2S U18491 ( .A(n29597), .B(n20376), .S(gray_img[1793]), .O(n18877) );
  ND2S U18492 ( .I1(n15884), .I2(n20568), .O(n20570) );
  MUX2S U18493 ( .A(n25928), .B(n20568), .S(gray_img[761]), .O(n20569) );
  AO12S U18494 ( .B1(n15931), .B2(n26841), .A1(n26723), .O(n14458) );
  MUX2S U18495 ( .A(n29587), .B(n20531), .S(gray_img[1673]), .O(n19538) );
  ND2S U18496 ( .I1(n28671), .I2(n28589), .O(n28592) );
  OA12S U18497 ( .B1(n29884), .B2(n28674), .A1(n28590), .O(n28591) );
  MUX2S U18498 ( .A(n15904), .B(n28672), .S(gray_img[545]), .O(n28590) );
  AO12S U18499 ( .B1(n15885), .B2(n26743), .A1(n26739), .O(n14450) );
  MUX2S U18500 ( .A(n27447), .B(n26741), .S(gray_img[337]), .O(n26739) );
  MUX2S U18501 ( .A(n25928), .B(n20452), .S(gray_img[889]), .O(n19520) );
  AO12S U18502 ( .B1(n15885), .B2(n28359), .A1(n28356), .O(n14361) );
  ND2S U18503 ( .I1(n15884), .I2(n20541), .O(n18481) );
  MUX2S U18504 ( .A(n29597), .B(n20541), .S(gray_img[1777]), .O(n18480) );
  MUX2S U18505 ( .A(n29597), .B(n20463), .S(gray_img[1641]), .O(n19534) );
  ND2S U18506 ( .I1(n15884), .I2(n20129), .O(n18621) );
  AO12S U18507 ( .B1(n15884), .B2(n28423), .A1(n28272), .O(n14394) );
  OA12S U18508 ( .B1(n25047), .B2(n25038), .A1(n25037), .O(n25039) );
  MUX2S U18509 ( .A(n25048), .B(n25047), .S(cnt_cro_y[1]), .O(n15747) );
  ND2S U18510 ( .I1(n15884), .I2(n20316), .O(n19767) );
  MUX2S U18511 ( .A(n29587), .B(n20316), .S(gray_img[1169]), .O(n19766) );
  MUX2S U18512 ( .A(n30050), .B(n23195), .S(gray_img[921]), .O(n23196) );
  MUX2S U18513 ( .A(n24958), .B(n24959), .S(cnt_cro_x[1]), .O(n15751) );
  MUX2S U18514 ( .A(n25928), .B(n20491), .S(gray_img[361]), .O(n19805) );
  AO12S U18515 ( .B1(n15931), .B2(n25653), .A1(n25650), .O(n14331) );
  ND2S U18516 ( .I1(n15932), .I2(n20684), .O(n20642) );
  MUX2S U18517 ( .A(n30050), .B(n20684), .S(gray_img[1473]), .O(n20641) );
  OA12S U18518 ( .B1(n29734), .B2(n23486), .A1(n23485), .O(n23487) );
  ND2S U18519 ( .I1(n26849), .I2(n23484), .O(n23488) );
  AO12S U18520 ( .B1(n24959), .B2(cnt_cro_x[2]), .A1(n24960), .O(n15750) );
  ND2S U18521 ( .I1(n30370), .I2(n30361), .O(n30363) );
  MUX2S U18522 ( .A(n24947), .B(n24946), .S(n24951), .O(n15761) );
  OR2S U18523 ( .I1(n30452), .I2(n19952), .O(n19954) );
  AN2S U18524 ( .I1(n30223), .I2(n30349), .O(gray_scale_2_n[7]) );
  AN2S U18525 ( .I1(C551_DATA2_6), .I2(n30349), .O(gray_scale_2_n[6]) );
  AN2S U18526 ( .I1(n30289), .I2(n30349), .O(gray_scale_1_n[9]) );
  AN2S U18527 ( .I1(n30286), .I2(n30349), .O(gray_scale_1_n[8]) );
  ND2S U18528 ( .I1(n30147), .I2(n30146), .O(n30149) );
  ND2S U18529 ( .I1(n30162), .I2(n30161), .O(n30164) );
  ND2S U18530 ( .I1(n30169), .I2(n30168), .O(n30172) );
  ND2S U18531 ( .I1(n30177), .I2(n30176), .O(n30178) );
  ND2S U18532 ( .I1(n30184), .I2(n30183), .O(n30185) );
  ND2S U18533 ( .I1(n30189), .I2(n30188), .O(n30191) );
  ND2S U18534 ( .I1(n30195), .I2(n30194), .O(n30196) );
  MUX2S U18535 ( .A(template_in_reg[7]), .B(template_reg[71]), .S(n30143), .O(
        n15661) );
  MUX2S U18536 ( .A(template_in_reg[6]), .B(template_reg[70]), .S(n30143), .O(
        n15662) );
  MUX2S U18537 ( .A(template_in_reg[5]), .B(template_reg[69]), .S(n30143), .O(
        n15663) );
  MUX2S U18538 ( .A(template_in_reg[4]), .B(template_reg[68]), .S(n30143), .O(
        n15664) );
  MUX2S U18539 ( .A(template_in_reg[3]), .B(template_reg[67]), .S(n30143), .O(
        n15665) );
  MUX2S U18540 ( .A(template_in_reg[2]), .B(template_reg[66]), .S(n30143), .O(
        n15666) );
  MUX2S U18541 ( .A(template_in_reg[1]), .B(template_reg[65]), .S(n30143), .O(
        n15667) );
  MUX2S U18542 ( .A(template_in_reg[0]), .B(template_reg[64]), .S(n30143), .O(
        n15668) );
  MUX2S U18543 ( .A(template_in_reg[7]), .B(template_reg[63]), .S(n30144), .O(
        n15669) );
  MUX2S U18544 ( .A(template_in_reg[6]), .B(template_reg[62]), .S(n30144), .O(
        n15670) );
  MUX2S U18545 ( .A(template_in_reg[5]), .B(template_reg[61]), .S(n30144), .O(
        n15671) );
  MUX2S U18546 ( .A(template_in_reg[4]), .B(template_reg[60]), .S(n30144), .O(
        n15672) );
  MUX2S U18547 ( .A(template_in_reg[3]), .B(template_reg[59]), .S(n30144), .O(
        n15673) );
  MUX2S U18548 ( .A(template_in_reg[2]), .B(template_reg[58]), .S(n30144), .O(
        n15674) );
  MUX2S U18549 ( .A(template_in_reg[1]), .B(template_reg[57]), .S(n30144), .O(
        n15675) );
  MUX2S U18550 ( .A(template_in_reg[0]), .B(template_reg[56]), .S(n30144), .O(
        n15676) );
  MUX2S U18551 ( .A(template_in_reg[7]), .B(template_reg[55]), .S(n30145), .O(
        n15677) );
  MUX2S U18552 ( .A(template_in_reg[6]), .B(template_reg[54]), .S(n30145), .O(
        n15678) );
  MUX2S U18553 ( .A(template_in_reg[5]), .B(template_reg[53]), .S(n30145), .O(
        n15679) );
  MUX2S U18554 ( .A(template_in_reg[4]), .B(template_reg[52]), .S(n30145), .O(
        n15680) );
  MUX2S U18555 ( .A(template_in_reg[3]), .B(template_reg[51]), .S(n30145), .O(
        n15681) );
  MUX2S U18556 ( .A(template_in_reg[2]), .B(template_reg[50]), .S(n30145), .O(
        n15682) );
  MUX2S U18557 ( .A(template_in_reg[1]), .B(template_reg[49]), .S(n30145), .O(
        n15683) );
  MUX2S U18558 ( .A(template_in_reg[0]), .B(template_reg[48]), .S(n30145), .O(
        n15684) );
  MUX2S U18559 ( .A(template_in_reg[7]), .B(template_reg[23]), .S(n30138), .O(
        n15709) );
  MUX2S U18560 ( .A(template_in_reg[6]), .B(template_reg[22]), .S(n30138), .O(
        n15710) );
  MUX2S U18561 ( .A(template_in_reg[5]), .B(template_reg[21]), .S(n30138), .O(
        n15711) );
  MUX2S U18562 ( .A(template_in_reg[4]), .B(template_reg[20]), .S(n30138), .O(
        n15712) );
  MUX2S U18563 ( .A(template_in_reg[3]), .B(template_reg[19]), .S(n30138), .O(
        n15713) );
  MUX2S U18564 ( .A(template_in_reg[2]), .B(template_reg[18]), .S(n30138), .O(
        n15714) );
  MUX2S U18565 ( .A(template_in_reg[1]), .B(template_reg[17]), .S(n30138), .O(
        n15715) );
  MUX2S U18566 ( .A(template_in_reg[0]), .B(template_reg[16]), .S(n30138), .O(
        n15716) );
  MUX2S U18567 ( .A(template_in_reg[7]), .B(template_reg[15]), .S(n30137), .O(
        n15717) );
  MUX2S U18568 ( .A(template_in_reg[6]), .B(template_reg[14]), .S(n30137), .O(
        n15718) );
  MUX2S U18569 ( .A(template_in_reg[5]), .B(template_reg[13]), .S(n30137), .O(
        n15719) );
  MUX2S U18570 ( .A(template_in_reg[4]), .B(template_reg[12]), .S(n30137), .O(
        n15720) );
  MUX2S U18571 ( .A(template_in_reg[3]), .B(template_reg[11]), .S(n30137), .O(
        n15721) );
  MUX2S U18572 ( .A(template_in_reg[2]), .B(template_reg[10]), .S(n30137), .O(
        n15722) );
  MUX2S U18573 ( .A(template_in_reg[1]), .B(template_reg[9]), .S(n30137), .O(
        n15723) );
  MUX2S U18574 ( .A(template_in_reg[0]), .B(template_reg[8]), .S(n30137), .O(
        n15724) );
  MUX2S U18575 ( .A(template_in_reg[7]), .B(template_reg[7]), .S(n30139), .O(
        n15725) );
  MUX2S U18576 ( .A(template_in_reg[6]), .B(template_reg[6]), .S(n30139), .O(
        n15726) );
  MUX2S U18577 ( .A(template_in_reg[5]), .B(template_reg[5]), .S(n30139), .O(
        n15727) );
  MUX2S U18578 ( .A(template_in_reg[4]), .B(template_reg[4]), .S(n30139), .O(
        n15728) );
  MUX2S U18579 ( .A(template_in_reg[3]), .B(template_reg[3]), .S(n30139), .O(
        n15729) );
  MUX2S U18580 ( .A(template_in_reg[2]), .B(template_reg[2]), .S(n30139), .O(
        n15730) );
  MUX2S U18581 ( .A(template_in_reg[1]), .B(template_reg[1]), .S(n30139), .O(
        n15731) );
  MUX2S U18582 ( .A(template_in_reg[0]), .B(template_reg[0]), .S(n30139), .O(
        n15732) );
  ND2S U18583 ( .I1(n20228), .I2(n20227), .O(n15469) );
  MUX2S U18584 ( .A(n29566), .B(n25942), .S(gray_img[2039]), .O(n20227) );
  ND2S U18585 ( .I1(n19974), .I2(n19973), .O(n15470) );
  MUX2S U18586 ( .A(n30005), .B(n20608), .S(gray_img[2031]), .O(n19973) );
  AO12S U18587 ( .B1(n15892), .B2(n25836), .A1(n25064), .O(n15471) );
  MUX2S U18588 ( .A(n25834), .B(n27447), .S(n25848), .O(n25064) );
  AO12S U18589 ( .B1(n15892), .B2(n25473), .A1(n24980), .O(n15472) );
  MUX2S U18590 ( .A(n25471), .B(n27447), .S(n24979), .O(n24980) );
  AO12S U18591 ( .B1(n15892), .B2(n25761), .A1(n24971), .O(n15473) );
  MUX2S U18592 ( .A(n27447), .B(n25759), .S(gray_img[2007]), .O(n24971) );
  AO12S U18593 ( .B1(n15892), .B2(n28803), .A1(n25002), .O(n15474) );
  MUX2S U18594 ( .A(n28801), .B(n15889), .S(n25001), .O(n25002) );
  ND2S U18595 ( .I1(n20211), .I2(n20210), .O(n15475) );
  MUX2S U18596 ( .A(n30044), .B(n20209), .S(gray_img[1991]), .O(n20211) );
  ND2S U18597 ( .I1(n20049), .I2(n20048), .O(n15476) );
  MUX2S U18598 ( .A(n29566), .B(n20746), .S(gray_img[1983]), .O(n20048) );
  ND2S U18599 ( .I1(n20208), .I2(n20207), .O(n15477) );
  MUX2S U18600 ( .A(n29597), .B(n20849), .S(gray_img[1975]), .O(n20208) );
  ND2S U18601 ( .I1(n20204), .I2(n20203), .O(n15478) );
  ND2S U18602 ( .I1(n20329), .I2(n20328), .O(n15479) );
  ND2S U18603 ( .I1(n19972), .I2(n19971), .O(n15480) );
  MUX2S U18604 ( .A(n20830), .B(n19970), .S(gray_img[1951]), .O(n19972) );
  ND2S U18605 ( .I1(n20220), .I2(n20219), .O(n15481) );
  MUX2S U18606 ( .A(n30050), .B(n20389), .S(gray_img[1943]), .O(n20220) );
  ND2S U18607 ( .I1(n20053), .I2(n20052), .O(n15482) );
  MUX2S U18608 ( .A(n30050), .B(n20424), .S(gray_img[1935]), .O(n20052) );
  ND2S U18609 ( .I1(n20226), .I2(n20225), .O(n15483) );
  MUX2S U18610 ( .A(n20842), .B(n20373), .S(gray_img[1927]), .O(n20226) );
  ND2S U18611 ( .I1(n20058), .I2(n20057), .O(n15484) );
  MUX2S U18612 ( .A(n29597), .B(n20430), .S(gray_img[1919]), .O(n20057) );
  ND2S U18613 ( .I1(n20065), .I2(n20064), .O(n15485) );
  MUX2S U18614 ( .A(n30044), .B(n20063), .S(gray_img[1911]), .O(n20064) );
  ND2S U18615 ( .I1(n20075), .I2(n20074), .O(n15486) );
  MUX2S U18616 ( .A(n30056), .B(n20544), .S(gray_img[1903]), .O(n20074) );
  ND2S U18617 ( .I1(n15889), .I2(n24975), .O(n24976) );
  AO12S U18618 ( .B1(n15892), .B2(n25460), .A1(n24969), .O(n15489) );
  ND2S U18619 ( .I1(n15889), .I2(n25004), .O(n25005) );
  ND2S U18620 ( .I1(n19967), .I2(n19966), .O(n15491) );
  MUX2S U18621 ( .A(n29566), .B(n20504), .S(gray_img[1863]), .O(n19966) );
  ND2S U18622 ( .I1(n20081), .I2(n20080), .O(n15492) );
  MUX2S U18623 ( .A(n29566), .B(n20740), .S(gray_img[1855]), .O(n20080) );
  ND2S U18624 ( .I1(n20175), .I2(n20174), .O(n15493) );
  MUX2S U18625 ( .A(n29597), .B(n20862), .S(gray_img[1847]), .O(n20175) );
  ND2S U18626 ( .I1(n20144), .I2(n20143), .O(n15494) );
  ND2S U18627 ( .I1(n20158), .I2(n20157), .O(n15495) );
  ND2S U18628 ( .I1(n20141), .I2(n20140), .O(n15496) );
  MUX2S U18629 ( .A(n29587), .B(n20296), .S(gray_img[1823]), .O(n20141) );
  ND2S U18630 ( .I1(n20341), .I2(n20340), .O(n15497) );
  MUX2S U18631 ( .A(n29597), .B(n20354), .S(gray_img[1815]), .O(n20341) );
  ND2S U18632 ( .I1(n20090), .I2(n20089), .O(n15498) );
  ND2S U18633 ( .I1(n20139), .I2(n20138), .O(n15499) );
  MUX2S U18634 ( .A(n29597), .B(n20376), .S(gray_img[1799]), .O(n20139) );
  ND2S U18635 ( .I1(n20034), .I2(n20033), .O(n15500) );
  MUX2S U18636 ( .A(n29597), .B(n20547), .S(gray_img[1791]), .O(n20033) );
  ND2S U18637 ( .I1(n20047), .I2(n20046), .O(n15501) );
  ND2S U18638 ( .I1(n19959), .I2(n19958), .O(n15502) );
  MUX2S U18639 ( .A(n30050), .B(n20449), .S(gray_img[1775]), .O(n19958) );
  AO12S U18640 ( .B1(n15892), .B2(n25778), .A1(n25060), .O(n15503) );
  MUX2S U18641 ( .A(n27447), .B(n25776), .S(gray_img[1767]), .O(n25060) );
  AO12S U18642 ( .B1(n15892), .B2(n25510), .A1(n24995), .O(n15504) );
  MUX2S U18643 ( .A(n27447), .B(n25508), .S(gray_img[1759]), .O(n24995) );
  AO12S U18644 ( .B1(n15892), .B2(n25498), .A1(n24991), .O(n15505) );
  MUX2S U18645 ( .A(n28534), .B(n25496), .S(gray_img[1751]), .O(n24991) );
  ND2S U18646 ( .I1(n19957), .I2(n19956), .O(n15507) );
  MUX2S U18647 ( .A(n29587), .B(n19955), .S(gray_img[1735]), .O(n19956) );
  ND2S U18648 ( .I1(n20092), .I2(n20091), .O(n15508) );
  MUX2S U18649 ( .A(n30056), .B(n20737), .S(gray_img[1727]), .O(n20091) );
  ND2S U18650 ( .I1(n20153), .I2(n20152), .O(n15509) );
  MUX2S U18651 ( .A(n30044), .B(n20846), .S(gray_img[1719]), .O(n20153) );
  ND2S U18652 ( .I1(n20188), .I2(n20187), .O(n15510) );
  MUX2S U18653 ( .A(n30056), .B(n20827), .S(gray_img[1711]), .O(n20188) );
  ND2S U18654 ( .I1(n20165), .I2(n20164), .O(n15511) );
  MUX2S U18655 ( .A(n30056), .B(n20787), .S(gray_img[1703]), .O(n20165) );
  ND2S U18656 ( .I1(n20199), .I2(n20198), .O(n15512) );
  MUX2S U18657 ( .A(n30056), .B(n20599), .S(gray_img[1695]), .O(n20199) );
  ND2S U18658 ( .I1(n20218), .I2(n20217), .O(n15513) );
  MUX2S U18659 ( .A(n29566), .B(n20605), .S(gray_img[1687]), .O(n20218) );
  ND2S U18660 ( .I1(n20028), .I2(n20027), .O(n15514) );
  MUX2S U18661 ( .A(n29587), .B(n20531), .S(gray_img[1679]), .O(n20027) );
  ND2S U18662 ( .I1(n20173), .I2(n20172), .O(n15515) );
  MUX2S U18663 ( .A(n29566), .B(n20583), .S(gray_img[1671]), .O(n20173) );
  ND2S U18664 ( .I1(n20069), .I2(n20068), .O(n15516) );
  ND2S U18665 ( .I1(n20107), .I2(n20106), .O(n15517) );
  ND2S U18666 ( .I1(n19963), .I2(n19962), .O(n15518) );
  MUX2S U18667 ( .A(n29597), .B(n20463), .S(gray_img[1647]), .O(n19962) );
  AO12S U18668 ( .B1(n15892), .B2(n25899), .A1(n25056), .O(n15519) );
  MUX2S U18669 ( .A(n15889), .B(n25897), .S(gray_img[1639]), .O(n25056) );
  AO12S U18670 ( .B1(n15892), .B2(n25576), .A1(n24993), .O(n15520) );
  MUX2S U18671 ( .A(n27447), .B(n25574), .S(gray_img[1631]), .O(n24993) );
  AO12S U18672 ( .B1(n15892), .B2(n25494), .A1(n24989), .O(n15521) );
  MUX2S U18673 ( .A(n27447), .B(n25492), .S(gray_img[1623]), .O(n24989) );
  ND2S U18674 ( .I1(n19965), .I2(n19964), .O(n15523) );
  MUX2S U18675 ( .A(n29566), .B(n20528), .S(gray_img[1607]), .O(n19964) );
  ND2S U18676 ( .I1(n20039), .I2(n20038), .O(n15524) );
  MUX2S U18677 ( .A(n30050), .B(n20731), .S(gray_img[1599]), .O(n20038) );
  ND2S U18678 ( .I1(n20171), .I2(n20170), .O(n15525) );
  MUX2S U18679 ( .A(n30056), .B(n20839), .S(gray_img[1591]), .O(n20171) );
  ND2S U18680 ( .I1(n20222), .I2(n20221), .O(n15526) );
  MUX2S U18681 ( .A(n30050), .B(n20395), .S(gray_img[1583]), .O(n20222) );
  ND2S U18682 ( .I1(n20216), .I2(n20215), .O(n15527) );
  MUX2S U18683 ( .A(n30056), .B(n20824), .S(gray_img[1575]), .O(n20216) );
  ND2S U18684 ( .I1(n19969), .I2(n19968), .O(n15528) );
  MUX2S U18685 ( .A(n29597), .B(n20596), .S(gray_img[1567]), .O(n19969) );
  ND2S U18686 ( .I1(n20224), .I2(n20223), .O(n15529) );
  MUX2S U18687 ( .A(n20830), .B(n20602), .S(gray_img[1559]), .O(n20224) );
  ND2S U18688 ( .I1(n19961), .I2(n19960), .O(n15530) );
  MUX2S U18689 ( .A(n29587), .B(n20550), .S(gray_img[1551]), .O(n19960) );
  ND2S U18690 ( .I1(n20876), .I2(n20875), .O(n15531) );
  MUX2S U18691 ( .A(n29597), .B(n20881), .S(gray_img[1543]), .O(n20876) );
  ND2S U18692 ( .I1(n20119), .I2(n20118), .O(n15532) );
  MUX2S U18693 ( .A(n30056), .B(n20556), .S(gray_img[1535]), .O(n20118) );
  ND2S U18694 ( .I1(n20105), .I2(n20104), .O(n15533) );
  ND2S U18695 ( .I1(n20086), .I2(n20085), .O(n15534) );
  MUX2S U18696 ( .A(n29566), .B(n20440), .S(gray_img[1519]), .O(n20085) );
  AO12S U18697 ( .B1(n15892), .B2(n27971), .A1(n25295), .O(n15535) );
  MUX2S U18698 ( .A(n28534), .B(n27969), .S(gray_img[1511]), .O(n25295) );
  AO12S U18699 ( .B1(n15892), .B2(n28355), .A1(n25184), .O(n15536) );
  MUX2S U18700 ( .A(n27447), .B(n28353), .S(gray_img[1503]), .O(n25184) );
  AO12S U18701 ( .B1(n15892), .B2(n28342), .A1(n25180), .O(n15537) );
  MUX2S U18702 ( .A(n15889), .B(n28340), .S(gray_img[1495]), .O(n25180) );
  ND2S U18703 ( .I1(n27447), .I2(n25199), .O(n25200) );
  ND2S U18704 ( .I1(n20067), .I2(n20066), .O(n15539) );
  MUX2S U18705 ( .A(n30050), .B(n20684), .S(gray_img[1479]), .O(n20066) );
  ND2S U18706 ( .I1(n20077), .I2(n20076), .O(n15540) );
  MUX2S U18707 ( .A(n30044), .B(n20709), .S(gray_img[1471]), .O(n20076) );
  ND2S U18708 ( .I1(n20181), .I2(n20180), .O(n15541) );
  MUX2S U18709 ( .A(n20830), .B(n20821), .S(gray_img[1463]), .O(n20181) );
  ND2S U18710 ( .I1(n20179), .I2(n20178), .O(n15542) );
  MUX2S U18711 ( .A(n20830), .B(n20814), .S(gray_img[1455]), .O(n20179) );
  ND2S U18712 ( .I1(n20177), .I2(n20176), .O(n15543) );
  MUX2S U18713 ( .A(n30050), .B(n20811), .S(gray_img[1447]), .O(n20177) );
  ND2S U18714 ( .I1(n20169), .I2(n20168), .O(n15544) );
  MUX2S U18715 ( .A(n30056), .B(n20293), .S(gray_img[1439]), .O(n20169) );
  ND2S U18716 ( .I1(n20195), .I2(n20194), .O(n15545) );
  MUX2S U18717 ( .A(n20842), .B(n20193), .S(gray_img[1431]), .O(n20195) );
  ND2S U18718 ( .I1(n20037), .I2(n20036), .O(n15546) );
  MUX2S U18719 ( .A(n29566), .B(n20035), .S(gray_img[1423]), .O(n20036) );
  ND2S U18720 ( .I1(n20190), .I2(n20189), .O(n15547) );
  ND2S U18721 ( .I1(n20113), .I2(n20112), .O(n15548) );
  MUX2S U18722 ( .A(n30044), .B(n20571), .S(gray_img[1407]), .O(n20112) );
  ND2S U18723 ( .I1(n20094), .I2(n20093), .O(n15549) );
  MUX2S U18724 ( .A(n30050), .B(n20517), .S(gray_img[1399]), .O(n20093) );
  ND2S U18725 ( .I1(n20096), .I2(n20095), .O(n15550) );
  MUX2S U18726 ( .A(n30050), .B(n20722), .S(gray_img[1391]), .O(n20095) );
  ND2S U18727 ( .I1(n15889), .I2(n28002), .O(n25289) );
  AO12S U18728 ( .B1(n25112), .B2(n28359), .A1(n25182), .O(n15552) );
  MUX2S U18729 ( .A(n27447), .B(n28357), .S(gray_img[1375]), .O(n25182) );
  AO12S U18730 ( .B1(n15892), .B2(n28596), .A1(n25178), .O(n15553) );
  MUX2S U18731 ( .A(n28534), .B(n28594), .S(gray_img[1367]), .O(n25178) );
  ND2S U18732 ( .I1(n15889), .I2(n25203), .O(n25204) );
  ND2S U18733 ( .I1(n20079), .I2(n20078), .O(n15555) );
  MUX2S U18734 ( .A(n29587), .B(n20734), .S(gray_img[1351]), .O(n20078) );
  ND2S U18735 ( .I1(n20032), .I2(n20031), .O(n15556) );
  ND2S U18736 ( .I1(n20137), .I2(n20136), .O(n15557) );
  MUX2S U18737 ( .A(n30050), .B(n20833), .S(gray_img[1335]), .O(n20137) );
  ND2S U18738 ( .I1(n20133), .I2(n20132), .O(n15558) );
  MUX2S U18739 ( .A(n29566), .B(n20836), .S(gray_img[1327]), .O(n20133) );
  ND2S U18740 ( .I1(n20151), .I2(n20150), .O(n15559) );
  MUX2S U18741 ( .A(n30050), .B(n20843), .S(gray_img[1319]), .O(n20151) );
  ND2S U18742 ( .I1(n20131), .I2(n20130), .O(n15560) );
  ND2S U18743 ( .I1(n20146), .I2(n20145), .O(n15561) );
  MUX2S U18744 ( .A(n29566), .B(n20362), .S(gray_img[1303]), .O(n20146) );
  ND2S U18745 ( .I1(n20041), .I2(n20040), .O(n15562) );
  ND2S U18746 ( .I1(n20135), .I2(n20134), .O(n15563) );
  MUX2S U18747 ( .A(n29587), .B(n20392), .S(gray_img[1287]), .O(n20135) );
  ND2S U18748 ( .I1(n20115), .I2(n20114), .O(n15564) );
  ND2S U18749 ( .I1(n20071), .I2(n20070), .O(n15565) );
  ND2S U18750 ( .I1(n20103), .I2(n20102), .O(n15566) );
  MUX2S U18751 ( .A(n30044), .B(n20719), .S(gray_img[1263]), .O(n20102) );
  AO12S U18752 ( .B1(n20271), .B2(n28031), .A1(n25299), .O(n15567) );
  MUX2S U18753 ( .A(n15889), .B(n28029), .S(gray_img[1255]), .O(n25299) );
  AO12S U18754 ( .B1(n25112), .B2(n28288), .A1(n25174), .O(n15568) );
  MUX2S U18755 ( .A(n28534), .B(n28286), .S(gray_img[1247]), .O(n25174) );
  AO12S U18756 ( .B1(n20271), .B2(n28271), .A1(n25172), .O(n15569) );
  MUX2S U18757 ( .A(n15889), .B(n28269), .S(gray_img[1239]), .O(n25172) );
  AO12S U18758 ( .B1(n15892), .B2(n28475), .A1(n25186), .O(n15570) );
  MUX2S U18759 ( .A(n27447), .B(n28473), .S(gray_img[1231]), .O(n25186) );
  ND2S U18760 ( .I1(n20111), .I2(n20110), .O(n15571) );
  MUX2S U18761 ( .A(n29587), .B(n20702), .S(gray_img[1223]), .O(n20110) );
  ND2S U18762 ( .I1(n20264), .I2(n20263), .O(n15572) );
  MUX2S U18763 ( .A(n30044), .B(n20757), .S(gray_img[1215]), .O(n20263) );
  ND2S U18764 ( .I1(n20155), .I2(n20154), .O(n15573) );
  MUX2S U18765 ( .A(n30044), .B(n20857), .S(gray_img[1207]), .O(n20155) );
  ND2S U18766 ( .I1(n20248), .I2(n20247), .O(n15574) );
  MUX2S U18767 ( .A(n29597), .B(n20435), .S(gray_img[1199]), .O(n20247) );
  ND2S U18768 ( .I1(n20163), .I2(n20162), .O(n15575) );
  MUX2S U18769 ( .A(n30056), .B(n20379), .S(gray_img[1191]), .O(n20163) );
  ND2S U18770 ( .I1(n20161), .I2(n20160), .O(n15576) );
  MUX2S U18771 ( .A(n29597), .B(n20159), .S(gray_img[1183]), .O(n20161) );
  ND2S U18772 ( .I1(n20239), .I2(n20238), .O(n15577) );
  MUX2S U18773 ( .A(n29597), .B(n20316), .S(gray_img[1175]), .O(n20238) );
  ND2S U18774 ( .I1(n20117), .I2(n20116), .O(n15578) );
  MUX2S U18775 ( .A(n29566), .B(n20553), .S(gray_img[1167]), .O(n20116) );
  ND2S U18776 ( .I1(n20242), .I2(n20241), .O(n15579) );
  MUX2S U18777 ( .A(n29566), .B(n20240), .S(gray_img[1159]), .O(n20241) );
  ND2S U18778 ( .I1(n20121), .I2(n20120), .O(n15580) );
  MUX2S U18779 ( .A(n30050), .B(n20716), .S(gray_img[1151]), .O(n20120) );
  ND2S U18780 ( .I1(n20126), .I2(n20125), .O(n15581) );
  ND2S U18781 ( .I1(n20128), .I2(n20127), .O(n15582) );
  MUX2S U18782 ( .A(n30056), .B(n20728), .S(gray_img[1135]), .O(n20127) );
  AO12S U18783 ( .B1(n15892), .B2(n28092), .A1(n25303), .O(n15583) );
  MUX2S U18784 ( .A(n27447), .B(n28090), .S(gray_img[1127]), .O(n25303) );
  AO12S U18785 ( .B1(n15892), .B2(n28284), .A1(n25176), .O(n15584) );
  MUX2S U18786 ( .A(n27447), .B(n28282), .S(gray_img[1119]), .O(n25176) );
  AO12S U18787 ( .B1(n25112), .B2(n28423), .A1(n25170), .O(n15585) );
  MUX2S U18788 ( .A(n15889), .B(n28421), .S(gray_img[1111]), .O(n25170) );
  AO12S U18789 ( .B1(n15892), .B2(n28480), .A1(n25188), .O(n15586) );
  MUX2S U18790 ( .A(n28534), .B(n28478), .S(gray_img[1103]), .O(n25188) );
  ND2S U18791 ( .I1(n20088), .I2(n20087), .O(n15587) );
  MUX2S U18792 ( .A(n30050), .B(n20743), .S(gray_img[1095]), .O(n20087) );
  ND2S U18793 ( .I1(n20268), .I2(n20267), .O(n15588) );
  MUX2S U18794 ( .A(n30056), .B(n20760), .S(gray_img[1087]), .O(n20267) );
  ND2S U18795 ( .I1(n20197), .I2(n20196), .O(n15589) );
  MUX2S U18796 ( .A(n30044), .B(n20854), .S(gray_img[1079]), .O(n20197) );
  ND2S U18797 ( .I1(n20230), .I2(n20229), .O(n15590) );
  MUX2S U18798 ( .A(n29587), .B(n20611), .S(gray_img[1071]), .O(n20229) );
  ND2S U18799 ( .I1(n20206), .I2(n20205), .O(n15591) );
  MUX2S U18800 ( .A(n29566), .B(n20368), .S(gray_img[1063]), .O(n20206) );
  ND2S U18801 ( .I1(n20186), .I2(n20185), .O(n15592) );
  MUX2S U18802 ( .A(n30056), .B(n20184), .S(gray_img[1055]), .O(n20186) );
  ND2S U18803 ( .I1(n20257), .I2(n20256), .O(n15593) );
  MUX2S U18804 ( .A(n30056), .B(n20255), .S(gray_img[1047]), .O(n20256) );
  ND2S U18805 ( .I1(n20237), .I2(n20236), .O(n15594) );
  MUX2S U18806 ( .A(n29597), .B(n20235), .S(gray_img[1039]), .O(n20236) );
  ND2S U18807 ( .I1(n20244), .I2(n20243), .O(n15595) );
  MUX2S U18808 ( .A(n29566), .B(n20311), .S(gray_img[1031]), .O(n20243) );
  ND2S U18809 ( .I1(n20101), .I2(n20100), .O(n15596) );
  MUX2S U18810 ( .A(n15904), .B(n20099), .S(gray_img[1023]), .O(n20100) );
  ND2S U18811 ( .I1(n20045), .I2(n20044), .O(n15597) );
  MUX2S U18812 ( .A(n20842), .B(n20562), .S(gray_img[1015]), .O(n20044) );
  ND2S U18813 ( .I1(n20192), .I2(n20191), .O(n15598) );
  MUX2S U18814 ( .A(n30005), .B(n20384), .S(gray_img[1007]), .O(n20192) );
  AO12S U18815 ( .B1(n15892), .B2(n27829), .A1(n25338), .O(n15599) );
  MUX2S U18816 ( .A(n27447), .B(n27827), .S(gray_img[999]), .O(n25338) );
  AO12S U18817 ( .B1(n15892), .B2(n27081), .A1(n25350), .O(n15600) );
  MUX2S U18818 ( .A(n27447), .B(n27079), .S(gray_img[991]), .O(n25350) );
  AO12S U18819 ( .B1(n15892), .B2(n27065), .A1(n25346), .O(n15601) );
  MUX2S U18820 ( .A(n15889), .B(n27063), .S(gray_img[983]), .O(n25346) );
  AO12S U18821 ( .B1(n15892), .B2(n27261), .A1(n25166), .O(n15602) );
  MUX2S U18822 ( .A(n27447), .B(n27259), .S(gray_img[975]), .O(n25166) );
  ND2S U18823 ( .I1(n20201), .I2(n20200), .O(n15603) );
  MUX2S U18824 ( .A(n29587), .B(n20580), .S(gray_img[967]), .O(n20201) );
  ND2S U18825 ( .I1(n20062), .I2(n20061), .O(n15604) );
  MUX2S U18826 ( .A(n30005), .B(n20452), .S(gray_img[895]), .O(n20061) );
  ND2S U18827 ( .I1(n20026), .I2(n20025), .O(n15605) );
  MUX2S U18828 ( .A(n30005), .B(n20559), .S(gray_img[887]), .O(n20025) );
  ND2S U18829 ( .I1(n20214), .I2(n20213), .O(n15606) );
  MUX2S U18830 ( .A(n30005), .B(n20212), .S(gray_img[879]), .O(n20214) );
  AO12S U18831 ( .B1(n20271), .B2(n26224), .A1(n25332), .O(n15607) );
  MUX2S U18832 ( .A(n27447), .B(n26222), .S(gray_img[871]), .O(n25332) );
  AO12S U18833 ( .B1(n15892), .B2(n30065), .A1(n25354), .O(n15608) );
  MUX2S U18834 ( .A(n27447), .B(n30063), .S(gray_img[863]), .O(n25354) );
  AO12S U18835 ( .B1(n15892), .B2(n27069), .A1(n25360), .O(n15609) );
  MUX2S U18836 ( .A(n15889), .B(n27067), .S(gray_img[855]), .O(n25360) );
  AO12S U18837 ( .B1(n15892), .B2(n27190), .A1(n25168), .O(n15610) );
  MUX2S U18838 ( .A(n27447), .B(n27188), .S(gray_img[847]), .O(n25168) );
  ND2S U18839 ( .I1(n20278), .I2(n20277), .O(n15611) );
  MUX2S U18840 ( .A(n29587), .B(n20634), .S(gray_img[839]), .O(n20277) );
  ND2S U18841 ( .I1(n20043), .I2(n20042), .O(n15612) );
  MUX2S U18842 ( .A(n30005), .B(n20568), .S(gray_img[767]), .O(n20042) );
  ND2S U18843 ( .I1(n20056), .I2(n20055), .O(n15613) );
  MUX2S U18844 ( .A(n30005), .B(n20054), .S(gray_img[759]), .O(n20055) );
  ND2S U18845 ( .I1(n20183), .I2(n20182), .O(n15614) );
  MUX2S U18846 ( .A(n30005), .B(n20365), .S(gray_img[751]), .O(n20183) );
  AO12S U18847 ( .B1(n20271), .B2(n26155), .A1(n25344), .O(n15615) );
  MUX2S U18848 ( .A(n27447), .B(n26153), .S(gray_img[743]), .O(n25344) );
  AO12S U18849 ( .B1(n15892), .B2(n26996), .A1(n25143), .O(n15616) );
  AO12S U18850 ( .B1(n15892), .B2(n27009), .A1(n25147), .O(n15617) );
  MUX2S U18851 ( .A(n27447), .B(n27007), .S(gray_img[727]), .O(n25147) );
  AO12S U18852 ( .B1(n15892), .B2(n27243), .A1(n25155), .O(n15618) );
  MUX2S U18853 ( .A(n27241), .B(n27447), .S(n27158), .O(n25155) );
  ND2S U18854 ( .I1(n20254), .I2(n20253), .O(n15619) );
  MUX2S U18855 ( .A(n29597), .B(n20623), .S(gray_img[711]), .O(n20253) );
  ND2S U18856 ( .I1(n20030), .I2(n20029), .O(n15620) );
  MUX2S U18857 ( .A(n30005), .B(n20565), .S(gray_img[639]), .O(n20029) );
  ND2S U18858 ( .I1(n20060), .I2(n20059), .O(n15621) );
  MUX2S U18859 ( .A(n30050), .B(n20534), .S(gray_img[631]), .O(n20059) );
  ND2S U18860 ( .I1(n20276), .I2(n20275), .O(n15622) );
  AO12S U18861 ( .B1(n15892), .B2(n26160), .A1(n25336), .O(n15623) );
  MUX2S U18862 ( .A(n15889), .B(n26158), .S(gray_img[615]), .O(n25336) );
  AO12S U18863 ( .B1(n15892), .B2(n27105), .A1(n25141), .O(n15624) );
  MUX2S U18864 ( .A(n27447), .B(n27103), .S(gray_img[607]), .O(n25141) );
  AO12S U18865 ( .B1(n15892), .B2(n27013), .A1(n25145), .O(n15625) );
  MUX2S U18866 ( .A(n27447), .B(n27011), .S(gray_img[599]), .O(n25145) );
  AO12S U18867 ( .B1(n15892), .B2(n27133), .A1(n25157), .O(n15626) );
  MUX2S U18868 ( .A(n27131), .B(n27447), .S(n25158), .O(n25157) );
  ND2S U18869 ( .I1(n20167), .I2(n20166), .O(n15627) );
  MUX2S U18870 ( .A(n29587), .B(n20591), .S(gray_img[583]), .O(n20167) );
  ND2S U18871 ( .I1(n20073), .I2(n20072), .O(n15628) );
  MUX2S U18872 ( .A(n30056), .B(n20472), .S(gray_img[511]), .O(n20072) );
  ND2S U18873 ( .I1(n20051), .I2(n20050), .O(n15629) );
  MUX2S U18874 ( .A(n30044), .B(n20477), .S(gray_img[503]), .O(n20050) );
  ND2S U18875 ( .I1(n20232), .I2(n20231), .O(n15630) );
  MUX2S U18876 ( .A(n29587), .B(n20480), .S(gray_img[495]), .O(n20231) );
  AO12S U18877 ( .B1(n15892), .B2(n27774), .A1(n25130), .O(n15631) );
  MUX2S U18878 ( .A(n27447), .B(n27772), .S(gray_img[487]), .O(n25130) );
  AO12S U18879 ( .B1(n15892), .B2(n27352), .A1(n25236), .O(n15632) );
  MUX2S U18880 ( .A(n27350), .B(n27447), .S(n26786), .O(n25236) );
  AO12S U18881 ( .B1(n15892), .B2(n26747), .A1(n25234), .O(n15633) );
  MUX2S U18882 ( .A(n27447), .B(n26745), .S(gray_img[471]), .O(n25234) );
  AO12S U18883 ( .B1(n15892), .B2(n26942), .A1(n25369), .O(n15634) );
  MUX2S U18884 ( .A(n28534), .B(n26940), .S(gray_img[463]), .O(n25369) );
  ND2S U18885 ( .I1(n20259), .I2(n20258), .O(n15635) );
  ND2S U18886 ( .I1(n20098), .I2(n20097), .O(n15636) );
  MUX2S U18887 ( .A(n15904), .B(n20486), .S(gray_img[383]), .O(n20097) );
  ND2S U18888 ( .I1(n20109), .I2(n20108), .O(n15637) );
  MUX2S U18889 ( .A(n30050), .B(n20522), .S(gray_img[375]), .O(n20108) );
  ND2S U18890 ( .I1(n20246), .I2(n20245), .O(n15638) );
  MUX2S U18891 ( .A(n29587), .B(n20491), .S(gray_img[367]), .O(n20245) );
  AO12S U18892 ( .B1(n20271), .B2(n27449), .A1(n25132), .O(n15639) );
  MUX2S U18893 ( .A(n27447), .B(n27446), .S(gray_img[359]), .O(n25132) );
  AO12S U18894 ( .B1(n15892), .B2(n26759), .A1(n25238), .O(n15640) );
  MUX2S U18895 ( .A(n26757), .B(n15889), .S(n25239), .O(n25238) );
  AO12S U18896 ( .B1(n15892), .B2(n26743), .A1(n25232), .O(n15641) );
  MUX2S U18897 ( .A(n15889), .B(n26741), .S(gray_img[343]), .O(n25232) );
  AO12S U18898 ( .B1(n15892), .B2(n26861), .A1(n25364), .O(n15642) );
  MUX2S U18899 ( .A(n27447), .B(n26859), .S(gray_img[335]), .O(n25364) );
  ND2S U18900 ( .I1(n20149), .I2(n20148), .O(n15643) );
  MUX2S U18901 ( .A(n30005), .B(n20147), .S(gray_img[327]), .O(n20149) );
  ND2S U18902 ( .I1(n20123), .I2(n20122), .O(n15644) );
  MUX2S U18903 ( .A(n29597), .B(n20496), .S(gray_img[255]), .O(n20122) );
  ND2S U18904 ( .I1(n20262), .I2(n20261), .O(n15645) );
  MUX2S U18905 ( .A(n29597), .B(n20260), .S(gray_img[247]), .O(n20261) );
  ND2S U18906 ( .I1(n20250), .I2(n20249), .O(n15646) );
  MUX2S U18907 ( .A(n20620), .B(n20830), .S(n27406), .O(n20249) );
  AO12S U18908 ( .B1(n25112), .B2(n27390), .A1(n25122), .O(n15647) );
  MUX2S U18909 ( .A(n15889), .B(n27388), .S(gray_img[231]), .O(n25122) );
  AO12S U18910 ( .B1(n25112), .B2(n26726), .A1(n25226), .O(n15648) );
  MUX2S U18911 ( .A(n27447), .B(n26724), .S(gray_img[223]), .O(n25226) );
  AO12S U18912 ( .B1(n15892), .B2(n26841), .A1(n25228), .O(n15649) );
  MUX2S U18913 ( .A(n27447), .B(n26839), .S(gray_img[215]), .O(n25228) );
  AO12S U18914 ( .B1(n20271), .B2(n26883), .A1(n25260), .O(n15650) );
  MUX2S U18915 ( .A(n15889), .B(n26881), .S(gray_img[207]), .O(n25260) );
  ND2S U18916 ( .I1(n20270), .I2(n20269), .O(n15651) );
  MUX2S U18917 ( .A(n20631), .B(n29566), .S(n23614), .O(n20269) );
  ND2S U18918 ( .I1(n20084), .I2(n20083), .O(n15652) );
  MUX2S U18919 ( .A(n29587), .B(n20082), .S(gray_img[127]), .O(n20083) );
  ND2S U18920 ( .I1(n20266), .I2(n20265), .O(n15653) );
  MUX2S U18921 ( .A(n30050), .B(n20499), .S(gray_img[119]), .O(n20265) );
  ND2S U18922 ( .I1(n20252), .I2(n20251), .O(n15654) );
  MUX2S U18923 ( .A(n20617), .B(n20830), .S(n25123), .O(n20251) );
  AO12S U18924 ( .B1(n15892), .B2(n27545), .A1(n25120), .O(n15655) );
  MUX2S U18925 ( .A(n27447), .B(n27543), .S(gray_img[103]), .O(n25120) );
  ND2S U18926 ( .I1(n15889), .I2(n25222), .O(n25223) );
  AO12S U18927 ( .B1(n15892), .B2(n26722), .A1(n25230), .O(n15657) );
  MUX2S U18928 ( .A(n28534), .B(n26720), .S(gray_img[87]), .O(n25230) );
  AO12S U18929 ( .B1(n25112), .B2(n26879), .A1(n25256), .O(n15658) );
  MUX2S U18930 ( .A(n27447), .B(n26877), .S(gray_img[79]), .O(n25256) );
  ND2S U18931 ( .I1(n20273), .I2(n20272), .O(n15659) );
  MUX2S U18932 ( .A(n20628), .B(n30005), .S(n23602), .O(n20272) );
  ND2S U18933 ( .I1(n20234), .I2(n20233), .O(n15660) );
  MUX2S U18934 ( .A(n29597), .B(n20614), .S(gray_img[2047]), .O(n20233) );
  ND2S U18935 ( .I1(n21988), .I2(n21987), .O(n15808) );
  AO12S U18936 ( .B1(n28847), .B2(n28819), .A1(n28818), .O(n13805) );
  ND2S U18937 ( .I1(n15888), .I2(n28840), .O(n28815) );
  ND2S U18938 ( .I1(n28727), .I2(n28726), .O(n28732) );
  OA12S U18939 ( .B1(n29734), .B2(n28730), .A1(n28729), .O(n28731) );
  AO12S U18940 ( .B1(n28724), .B2(n28723), .A1(n28722), .O(n13707) );
  MUX2S U18941 ( .A(n15904), .B(n28718), .S(gray_img[952]), .O(n28720) );
  AO12S U18942 ( .B1(n26096), .B2(n26095), .A1(n26094), .O(n13708) );
  MUX2S U18943 ( .A(n15904), .B(n26090), .S(gray_img[944]), .O(n26092) );
  ND2S U18944 ( .I1(n28806), .I2(n28805), .O(n28811) );
  MUX2S U18945 ( .A(n29566), .B(n28807), .S(gray_img[400]), .O(n28808) );
  AO12S U18946 ( .B1(n25619), .B2(n23293), .A1(n23292), .O(n13709) );
  MUX2S U18947 ( .A(n30044), .B(n25612), .S(gray_img[936]), .O(n23290) );
  OA12S U18948 ( .B1(n29734), .B2(n23586), .A1(n23585), .O(n23587) );
  ND2S U18949 ( .I1(n25758), .I2(n23583), .O(n23588) );
  OA12S U18950 ( .B1(n29734), .B2(n23363), .A1(n23362), .O(n23364) );
  ND2S U18951 ( .I1(n30128), .I2(n23361), .O(n23365) );
  AO12S U18952 ( .B1(n30038), .B2(n30037), .A1(n30036), .O(n13777) );
  ND3S U18953 ( .I1(n30035), .I2(n30034), .I3(n30033), .O(n30036) );
  MUX2S U18954 ( .A(n30050), .B(n30032), .S(gray_img[392]), .O(n30034) );
  ND2S U18955 ( .I1(n30020), .I2(n30019), .O(n30025) );
  OA12S U18956 ( .B1(n29734), .B2(n30023), .A1(n30022), .O(n30024) );
  AO12S U18957 ( .B1(n30109), .B2(n30108), .A1(n30107), .O(n13778) );
  MUX2S U18958 ( .A(n15904), .B(n30103), .S(gray_img[384]), .O(n30105) );
  AO12S U18959 ( .B1(n29604), .B2(n29603), .A1(n29602), .O(n13713) );
  MUX2S U18960 ( .A(n29597), .B(n29598), .S(gray_img[904]), .O(n29600) );
  AO12S U18961 ( .B1(n30098), .B2(n30097), .A1(n30096), .O(n13714) );
  MUX2S U18962 ( .A(n30044), .B(n30092), .S(gray_img[896]), .O(n30094) );
  AO12S U18963 ( .B1(n26080), .B2(n26052), .A1(n26051), .O(n13715) );
  MUX2S U18964 ( .A(n15904), .B(n26073), .S(gray_img[824]), .O(n26049) );
  AO12S U18965 ( .B1(n25936), .B2(n25907), .A1(n25906), .O(n13716) );
  ND3S U18966 ( .I1(n25905), .I2(n25904), .I3(n25903), .O(n25906) );
  MUX2S U18967 ( .A(n25928), .B(n25929), .S(gray_img[816]), .O(n25904) );
  AO12S U18968 ( .B1(n25750), .B2(n25749), .A1(n25748), .O(n13718) );
  MUX2S U18969 ( .A(n25928), .B(n25744), .S(gray_img[800]), .O(n25746) );
  AO12S U18970 ( .B1(n29273), .B2(n29265), .A1(n29264), .O(n13719) );
  MUX2S U18971 ( .A(n29566), .B(n29266), .S(gray_img[792]), .O(n29262) );
  AO12S U18972 ( .B1(n29192), .B2(n29191), .A1(n29190), .O(n13720) );
  MUX2S U18973 ( .A(n15904), .B(n29186), .S(gray_img[784]), .O(n29188) );
  AO12S U18974 ( .B1(n29487), .B2(n29486), .A1(n29485), .O(n13722) );
  ND3S U18975 ( .I1(n29484), .I2(n29483), .I3(n29482), .O(n29485) );
  ND2S U18976 ( .I1(n28247), .I2(n28216), .O(n28219) );
  OA12S U18977 ( .B1(n29734), .B2(n28250), .A1(n28217), .O(n28218) );
  ND2S U18978 ( .I1(n28136), .I2(n28135), .O(n28141) );
  OA12S U18979 ( .B1(n29734), .B2(n28139), .A1(n28138), .O(n28140) );
  AO12S U18980 ( .B1(n28214), .B2(n28213), .A1(n28212), .O(n13724) );
  MUX2S U18981 ( .A(n30005), .B(n28208), .S(gray_img[688]), .O(n28210) );
  OA12S U18982 ( .B1(n29734), .B2(n28709), .A1(n28681), .O(n28682) );
  AO12S U18983 ( .B1(n28607), .B2(n28606), .A1(n28605), .O(n13725) );
  ND3S U18984 ( .I1(n28604), .I2(n28603), .I3(n28602), .O(n28605) );
  MUX2S U18985 ( .A(n15904), .B(n28601), .S(gray_img[680]), .O(n28603) );
  AO12S U18986 ( .B1(n29381), .B2(n29358), .A1(n29357), .O(n14267) );
  MUX2S U18987 ( .A(n29566), .B(n29374), .S(gray_img[264]), .O(n29355) );
  AO12S U18988 ( .B1(n29350), .B2(n29349), .A1(n29348), .O(n13727) );
  MUX2S U18989 ( .A(n29587), .B(n29344), .S(gray_img[664]), .O(n29346) );
  AO12S U18990 ( .B1(n29904), .B2(n29903), .A1(n29902), .O(n13737) );
  MUX2S U18991 ( .A(n15904), .B(n29898), .S(gray_img[648]), .O(n29900) );
  ND2S U18992 ( .I1(n29993), .I2(n29992), .O(n29998) );
  OA12S U18993 ( .B1(n29734), .B2(n29996), .A1(n29995), .O(n29997) );
  AO12S U18994 ( .B1(n28128), .B2(n28100), .A1(n28099), .O(n13740) );
  MUX2S U18995 ( .A(n30056), .B(n28121), .S(gray_img[560]), .O(n28097) );
  ND2S U18996 ( .I1(n28671), .I2(n28670), .O(n28676) );
  OA12S U18997 ( .B1(n29734), .B2(n28674), .A1(n28673), .O(n28675) );
  AO12S U18998 ( .B1(n28950), .B2(n28942), .A1(n28941), .O(n13743) );
  ND2S U18999 ( .I1(n29043), .I2(n29042), .O(n29048) );
  MUX2S U19000 ( .A(n29597), .B(n29044), .S(gray_img[528]), .O(n29045) );
  OA12S U19001 ( .B1(n29734), .B2(n29883), .A1(n29855), .O(n29856) );
  MUX2S U19002 ( .A(n30005), .B(n29881), .S(gray_img[520]), .O(n29855) );
  AO12S U19003 ( .B1(n30087), .B2(n30086), .A1(n30085), .O(n13754) );
  MUX2S U19004 ( .A(n15904), .B(n30081), .S(gray_img[8]), .O(n30083) );
  AO12S U19005 ( .B1(n27851), .B2(n27850), .A1(n27849), .O(n13762) );
  AO12S U19006 ( .B1(n27840), .B2(n27839), .A1(n27838), .O(n13764) );
  MUX2S U19007 ( .A(n15904), .B(n27834), .S(gray_img[432]), .O(n27836) );
  AO12S U19008 ( .B1(n30076), .B2(n30075), .A1(n30074), .O(n13772) );
  MUX2S U19009 ( .A(n30044), .B(n30070), .S(gray_img[144]), .O(n30072) );
  ND2S U19010 ( .I1(n23121), .I2(n23089), .O(n23093) );
  OA12S U19011 ( .B1(n29734), .B2(n27224), .A1(n23294), .O(n23298) );
  ND2S U19012 ( .I1(n27226), .I2(n23296), .O(n23297) );
  MUX2S U19013 ( .A(n30044), .B(n27222), .S(gray_img[416]), .O(n23294) );
  AO12S U19014 ( .B1(n26489), .B2(n26488), .A1(n26487), .O(n13779) );
  MUX2S U19015 ( .A(n29587), .B(n26483), .S(gray_img[312]), .O(n26485) );
  OA12S U19016 ( .B1(n29734), .B2(n27254), .A1(n27246), .O(n27247) );
  ND2S U19017 ( .I1(n27251), .I2(n27245), .O(n27248) );
  MUX2S U19018 ( .A(n29597), .B(n27252), .S(gray_img[288]), .O(n27246) );
  AO12S U19019 ( .B1(n27821), .B2(n27793), .A1(n27792), .O(n13792) );
  MUX2S U19020 ( .A(n30005), .B(n27814), .S(gray_img[24]), .O(n27790) );
  AO12S U19021 ( .B1(n27785), .B2(n27784), .A1(n27783), .O(n13794) );
  MUX2S U19022 ( .A(n29597), .B(n27779), .S(gray_img[176]), .O(n27781) );
  OA12S U19023 ( .B1(n29734), .B2(n23414), .A1(n23413), .O(n23415) );
  ND2S U19024 ( .I1(n26939), .I2(n23411), .O(n23416) );
  AO12S U19025 ( .B1(n27708), .B2(n27707), .A1(n27706), .O(n13807) );
  AO12S U19026 ( .B1(n27556), .B2(n27555), .A1(n27554), .O(n13808) );
  OA12S U19027 ( .B1(n29734), .B2(n23628), .A1(n23627), .O(n23629) );
  ND2S U19028 ( .I1(n26931), .I2(n23625), .O(n23630) );
  MUX2S U19029 ( .A(n15889), .B(n25834), .S(gray_img[2016]), .O(n25835) );
  MUX2S U19030 ( .A(n27447), .B(n25471), .S(gray_img[2008]), .O(n25466) );
  MUX2S U19031 ( .A(n27447), .B(n25759), .S(gray_img[2000]), .O(n25760) );
  MUX2S U19032 ( .A(n15889), .B(n28801), .S(gray_img[1992]), .O(n28802) );
  MUX2S U19033 ( .A(n29566), .B(n20746), .S(gray_img[1976]), .O(n19116) );
  MUX2S U19034 ( .A(n29597), .B(n20849), .S(gray_img[1968]), .O(n19122) );
  MUX2S U19035 ( .A(n30044), .B(n19970), .S(gray_img[1944]), .O(n19344) );
  MUX2S U19036 ( .A(n29566), .B(n20389), .S(gray_img[1936]), .O(n19340) );
  MUX2S U19037 ( .A(n20842), .B(n20424), .S(gray_img[1928]), .O(n19334) );
  MUX2S U19038 ( .A(n20830), .B(n20373), .S(gray_img[1920]), .O(n19106) );
  MUX2S U19039 ( .A(n30050), .B(n20544), .S(gray_img[1896]), .O(n19028) );
  MUX2S U19040 ( .A(n15889), .B(n25475), .S(gray_img[1880]), .O(n25476) );
  MUX2S U19041 ( .A(n15889), .B(n25458), .S(gray_img[1872]), .O(n25454) );
  MUX2S U19042 ( .A(n15889), .B(n25629), .S(gray_img[1864]), .O(n25624) );
  MUX2S U19043 ( .A(n29587), .B(n20504), .S(gray_img[1856]), .O(n18979) );
  MUX2S U19044 ( .A(n29597), .B(n20740), .S(gray_img[1848]), .O(n19336) );
  MUX2S U19045 ( .A(n29597), .B(n20142), .S(gray_img[1832]), .O(n19040) );
  MUX2S U19046 ( .A(n29597), .B(n20354), .S(gray_img[1808]), .O(n20353) );
  MUX2S U19047 ( .A(n20808), .B(n20319), .S(gray_img[1800]), .O(n19342) );
  MUX2S U19048 ( .A(n29566), .B(n20376), .S(gray_img[1792]), .O(n19138) );
  MUX2S U19049 ( .A(n30050), .B(n20547), .S(gray_img[1784]), .O(n19083) );
  MUX2S U19050 ( .A(n29597), .B(n20541), .S(gray_img[1776]), .O(n19022) );
  MUX2S U19051 ( .A(n30056), .B(n20449), .S(gray_img[1768]), .O(n19156) );
  MUX2S U19052 ( .A(n15889), .B(n25508), .S(gray_img[1752]), .O(n25503) );
  MUX2S U19053 ( .A(n27447), .B(n25647), .S(gray_img[1736]), .O(n25642) );
  MUX2S U19054 ( .A(n29566), .B(n19955), .S(gray_img[1728]), .O(n19026) );
  MUX2S U19055 ( .A(n30050), .B(n20737), .S(gray_img[1720]), .O(n19104) );
  MUX2S U19056 ( .A(n20830), .B(n20846), .S(gray_img[1712]), .O(n19328) );
  MUX2S U19057 ( .A(n30050), .B(n20827), .S(gray_img[1704]), .O(n19118) );
  MUX2S U19058 ( .A(n30056), .B(n20787), .S(gray_img[1696]), .O(n19120) );
  MUX2S U19059 ( .A(n29597), .B(n20599), .S(gray_img[1688]), .O(n19034) );
  MUX2S U19060 ( .A(n29566), .B(n20531), .S(gray_img[1672]), .O(n19168) );
  MUX2S U19061 ( .A(n29587), .B(n20583), .S(gray_img[1664]), .O(n19020) );
  MUX2S U19062 ( .A(n29587), .B(n20525), .S(gray_img[1648]), .O(n19010) );
  MUX2S U19063 ( .A(n30050), .B(n20463), .S(gray_img[1640]), .O(n19136) );
  MUX2S U19064 ( .A(n15889), .B(n25897), .S(gray_img[1632]), .O(n25898) );
  MUX2S U19065 ( .A(n27447), .B(n25574), .S(gray_img[1624]), .O(n25575) );
  MUX2S U19066 ( .A(n27447), .B(n25651), .S(gray_img[1608]), .O(n25652) );
  MUX2S U19067 ( .A(n29587), .B(n20528), .S(gray_img[1600]), .O(n19166) );
  MUX2S U19068 ( .A(n30050), .B(n20731), .S(gray_img[1592]), .O(n19326) );
  MUX2S U19069 ( .A(n20830), .B(n20839), .S(gray_img[1584]), .O(n19102) );
  MUX2S U19070 ( .A(n30050), .B(n20395), .S(gray_img[1576]), .O(n19316) );
  MUX2S U19071 ( .A(n30056), .B(n20824), .S(gray_img[1568]), .O(n19322) );
  MUX2S U19072 ( .A(n30050), .B(n20550), .S(gray_img[1544]), .O(n19160) );
  MUX2S U19073 ( .A(n29566), .B(n20881), .S(gray_img[1536]), .O(n20883) );
  MUX2S U19074 ( .A(n30050), .B(n20556), .S(gray_img[1528]), .O(n18737) );
  MUX2S U19075 ( .A(n20842), .B(n20512), .S(gray_img[1520]), .O(n19012) );
  MUX2S U19076 ( .A(n30044), .B(n20440), .S(gray_img[1512]), .O(n19162) );
  AO12S U19077 ( .B1(n19092), .B2(n28342), .A1(n28335), .O(n13943) );
  MUX2S U19078 ( .A(n27447), .B(n28340), .S(gray_img[1488]), .O(n28335) );
  MUX2S U19079 ( .A(n20830), .B(n20709), .S(gray_img[1464]), .O(n19126) );
  MUX2S U19080 ( .A(n30044), .B(n20821), .S(gray_img[1456]), .O(n19036) );
  MUX2S U19081 ( .A(n29566), .B(n20814), .S(gray_img[1448]), .O(n19124) );
  MUX2S U19082 ( .A(n30056), .B(n20293), .S(gray_img[1432]), .O(n19094) );
  MUX2S U19083 ( .A(n20842), .B(n20193), .S(gray_img[1424]), .O(n19314) );
  MUX2S U19084 ( .A(n20842), .B(n20035), .S(gray_img[1416]), .O(n19324) );
  MUX2S U19085 ( .A(n30050), .B(n20571), .S(gray_img[1400]), .O(n19085) );
  MUX2S U19086 ( .A(n20808), .B(n20517), .S(gray_img[1392]), .O(n19144) );
  MUX2S U19087 ( .A(n20842), .B(n20722), .S(gray_img[1384]), .O(n19060) );
  AO12S U19088 ( .B1(n19092), .B2(n28203), .A1(n28202), .O(n13990) );
  MUX2S U19089 ( .A(n28534), .B(n28201), .S(gray_img[1376]), .O(n28202) );
  MUX2S U19090 ( .A(n29587), .B(n20734), .S(gray_img[1344]), .O(n19042) );
  MUX2S U19091 ( .A(n30056), .B(n20695), .S(gray_img[1336]), .O(n19080) );
  MUX2S U19092 ( .A(n30050), .B(n20833), .S(gray_img[1328]), .O(n19074) );
  MUX2S U19093 ( .A(n20842), .B(n20427), .S(gray_img[1288]), .O(n19142) );
  MUX2S U19094 ( .A(n30044), .B(n20655), .S(gray_img[1272]), .O(n18769) );
  MUX2S U19095 ( .A(n20808), .B(n20725), .S(gray_img[1264]), .O(n19150) );
  MUX2S U19096 ( .A(n30050), .B(n20702), .S(gray_img[1216]), .O(n19054) );
  ND2S U19097 ( .I1(n19739), .I2(n19738), .O(n14046) );
  MUX2S U19098 ( .A(n30056), .B(n20757), .S(gray_img[1208]), .O(n19738) );
  MUX2S U19099 ( .A(n30044), .B(n20857), .S(gray_img[1200]), .O(n19312) );
  MUX2S U19100 ( .A(n30044), .B(n20435), .S(gray_img[1192]), .O(n19674) );
  MUX2S U19101 ( .A(n29587), .B(n20379), .S(gray_img[1184]), .O(n19058) );
  MUX2S U19102 ( .A(n29597), .B(n20159), .S(gray_img[1176]), .O(n19100) );
  MUX2S U19103 ( .A(n15904), .B(n20316), .S(gray_img[1168]), .O(n19764) );
  MUX2S U19104 ( .A(n29587), .B(n20240), .S(gray_img[1152]), .O(n19708) );
  MUX2S U19105 ( .A(n20808), .B(n20124), .S(gray_img[1136]), .O(n19062) );
  MUX2S U19106 ( .A(n30056), .B(n20728), .S(gray_img[1128]), .O(n19066) );
  MUX2S U19107 ( .A(n27447), .B(n28090), .S(gray_img[1120]), .O(n28091) );
  MUX2S U19108 ( .A(n15889), .B(n28282), .S(gray_img[1112]), .O(n28283) );
  MUX2S U19109 ( .A(n30044), .B(n20854), .S(gray_img[1072]), .O(n19098) );
  MUX2S U19110 ( .A(n29597), .B(n20368), .S(gray_img[1056]), .O(n19064) );
  MUX2S U19111 ( .A(n29597), .B(n20235), .S(gray_img[1032]), .O(n19424) );
  MUX2S U19112 ( .A(n27447), .B(n27827), .S(gray_img[992]), .O(n27828) );
  MUX2S U19113 ( .A(n30005), .B(n20212), .S(gray_img[872]), .O(n19078) );
  ND2S U19114 ( .I1(n19927), .I2(n19926), .O(n14134) );
  MUX2S U19115 ( .A(n20634), .B(n30056), .S(n22990), .O(n19926) );
  MUX2S U19116 ( .A(n25928), .B(n20568), .S(gray_img[760]), .O(n19052) );
  ND2S U19117 ( .I1(n19880), .I2(n19879), .O(n14170) );
  MUX2S U19118 ( .A(n29032), .B(n20623), .S(gray_img[704]), .O(n19879) );
  MUX2S U19119 ( .A(n20842), .B(n20534), .S(gray_img[624]), .O(n19072) );
  ND2S U19120 ( .I1(n19860), .I2(n19859), .O(n14173) );
  MUX2S U19121 ( .A(n15904), .B(n20274), .S(gray_img[616]), .O(n19859) );
  MUX2S U19122 ( .A(n15889), .B(n27103), .S(gray_img[600]), .O(n27104) );
  MUX2S U19123 ( .A(n29587), .B(n20591), .S(gray_img[576]), .O(n19154) );
  MUX2S U19124 ( .A(n30050), .B(n20472), .S(gray_img[504]), .O(n19056) );
  MUX2S U19125 ( .A(n20808), .B(n20477), .S(gray_img[496]), .O(n19050) );
  MUX2S U19126 ( .A(n27447), .B(n27772), .S(gray_img[480]), .O(n27773) );
  AO12S U19127 ( .B1(n19092), .B2(n27352), .A1(n27351), .O(n14204) );
  MUX2S U19128 ( .A(n28534), .B(n27350), .S(gray_img[472]), .O(n27351) );
  MUX2S U19129 ( .A(n15889), .B(n26940), .S(gray_img[456]), .O(n26941) );
  ND2S U19130 ( .I1(n19886), .I2(n19885), .O(n14214) );
  MUX2S U19131 ( .A(n30050), .B(n20486), .S(gray_img[376]), .O(n19018) );
  MUX2S U19132 ( .A(n30044), .B(n20522), .S(gray_img[368]), .O(n19016) );
  MUX2S U19133 ( .A(n29597), .B(n20491), .S(gray_img[360]), .O(n19814) );
  MUX2S U19134 ( .A(n29566), .B(n20496), .S(gray_img[248]), .O(n19038) );
  ND2S U19135 ( .I1(n19747), .I2(n19746), .O(n14231) );
  MUX2S U19136 ( .A(n30050), .B(n20260), .S(gray_img[240]), .O(n19746) );
  MUX2S U19137 ( .A(n29597), .B(n20620), .S(gray_img[232]), .O(n19853) );
  MUX2S U19138 ( .A(n27447), .B(n27388), .S(gray_img[224]), .O(n27383) );
  ND2S U19139 ( .I1(n19901), .I2(n19900), .O(n14258) );
  MUX2S U19140 ( .A(n30044), .B(n20631), .S(gray_img[192]), .O(n19900) );
  MUX2S U19141 ( .A(n29597), .B(n20082), .S(gray_img[120]), .O(n19014) );
  MUX2S U19142 ( .A(n29566), .B(n20617), .S(gray_img[104]), .O(n19863) );
  MUX2S U19143 ( .A(n27447), .B(n27543), .S(gray_img[96]), .O(n27544) );
  OA222S U19144 ( .A1(n24868), .A2(n24867), .B1(n24866), .B2(n24865), .C1(
        n24864), .C2(n24863), .O(n24872) );
  ND2S U19145 ( .I1(n22217), .I2(n22216), .O(n15815) );
  AO12S U19146 ( .B1(n30120), .B2(n30119), .A1(n30118), .O(n13811) );
  MUX2S U19147 ( .A(n30005), .B(n30114), .S(gray_img[0]), .O(n30115) );
  AO12S U19148 ( .B1(n28847), .B2(n28846), .A1(n28845), .O(n14274) );
  ND2S U19149 ( .I1(n15932), .I2(n28840), .O(n28841) );
  MUX2S U19150 ( .A(n15904), .B(n28840), .S(gray_img[137]), .O(n28842) );
  AO12S U19151 ( .B1(n28724), .B2(n26085), .A1(n26084), .O(n13680) );
  ND2S U19152 ( .I1(n15932), .I2(n28718), .O(n26081) );
  MUX2S U19153 ( .A(n15904), .B(n28718), .S(gray_img[953]), .O(n26082) );
  AO12S U19154 ( .B1(n26096), .B2(n25941), .A1(n25940), .O(n13681) );
  ND2S U19155 ( .I1(n15928), .I2(n26090), .O(n25937) );
  MUX2S U19156 ( .A(n15904), .B(n26090), .S(gray_img[945]), .O(n25938) );
  AO12S U19157 ( .B1(n25758), .B2(n25757), .A1(n25756), .O(n13683) );
  ND2S U19158 ( .I1(n15932), .I2(n25751), .O(n25752) );
  MUX2S U19159 ( .A(n29566), .B(n25751), .S(gray_img[929]), .O(n25753) );
  AO12S U19160 ( .B1(n30128), .B2(n30127), .A1(n30126), .O(n14275) );
  ND2S U19161 ( .I1(n15932), .I2(n30121), .O(n30122) );
  MUX2S U19162 ( .A(n30044), .B(n30121), .S(gray_img[129]), .O(n30123) );
  AO12S U19163 ( .B1(n26080), .B2(n26079), .A1(n26078), .O(n13688) );
  ND2S U19164 ( .I1(n15932), .I2(n26073), .O(n26074) );
  MUX2S U19165 ( .A(n15904), .B(n26073), .S(gray_img[825]), .O(n26075) );
  AO12S U19166 ( .B1(n25936), .B2(n25935), .A1(n25934), .O(n13689) );
  MUX2S U19167 ( .A(n25928), .B(n25929), .S(gray_img[817]), .O(n25931) );
  OA12S U19168 ( .B1(n29884), .B2(n25607), .A1(n25606), .O(n25608) );
  MUX2S U19169 ( .A(n25928), .B(n25605), .S(gray_img[809]), .O(n25606) );
  AO12S U19170 ( .B1(n25750), .B2(n25719), .A1(n25718), .O(n13691) );
  ND2S U19171 ( .I1(n15929), .I2(n25744), .O(n25715) );
  MUX2S U19172 ( .A(n25928), .B(n25744), .S(gray_img[801]), .O(n25716) );
  AO12S U19173 ( .B1(n29273), .B2(n29272), .A1(n29271), .O(n13692) );
  ND2S U19174 ( .I1(n15932), .I2(n29266), .O(n29267) );
  MUX2S U19175 ( .A(n30050), .B(n29266), .S(gray_img[793]), .O(n29268) );
  AO12S U19176 ( .B1(n29192), .B2(n29161), .A1(n29160), .O(n13693) );
  ND2S U19177 ( .I1(n15932), .I2(n29186), .O(n29157) );
  MUX2S U19178 ( .A(n29597), .B(n29186), .S(gray_img[785]), .O(n29158) );
  AO12S U19179 ( .B1(n29487), .B2(n29456), .A1(n29455), .O(n13695) );
  MUX2S U19180 ( .A(n30056), .B(n29481), .S(gray_img[769]), .O(n29453) );
  ND2S U19181 ( .I1(n28247), .I2(n28236), .O(n28239) );
  OA12S U19182 ( .B1(n29884), .B2(n28250), .A1(n28237), .O(n28238) );
  MUX2S U19183 ( .A(n15904), .B(n28248), .S(gray_img[281]), .O(n28237) );
  ND2S U19184 ( .I1(n28136), .I2(n27954), .O(n27957) );
  OA12S U19185 ( .B1(n29884), .B2(n28139), .A1(n27955), .O(n27956) );
  MUX2S U19186 ( .A(n30005), .B(n28137), .S(gray_img[697]), .O(n27955) );
  AO12S U19187 ( .B1(n28607), .B2(n28464), .A1(n28463), .O(n13698) );
  ND2S U19188 ( .I1(n15932), .I2(n28601), .O(n28460) );
  MUX2S U19189 ( .A(n15904), .B(n28601), .S(gray_img[681]), .O(n28461) );
  AO12S U19190 ( .B1(n29381), .B2(n29380), .A1(n29379), .O(n13706) );
  ND2S U19191 ( .I1(n15932), .I2(n29374), .O(n29375) );
  MUX2S U19192 ( .A(n29587), .B(n29374), .S(gray_img[265]), .O(n29376) );
  AO12S U19193 ( .B1(n30087), .B2(n28852), .A1(n28851), .O(n13753) );
  ND2S U19194 ( .I1(n15932), .I2(n30081), .O(n28848) );
  MUX2S U19195 ( .A(n29587), .B(n30081), .S(gray_img[9]), .O(n28849) );
  AO12S U19196 ( .B1(n27851), .B2(n27826), .A1(n27825), .O(n13761) );
  MUX2S U19197 ( .A(n15904), .B(n27845), .S(gray_img[153]), .O(n27823) );
  AO12S U19198 ( .B1(n30076), .B2(n27329), .A1(n27328), .O(n13771) );
  ND2S U19199 ( .I1(n15932), .I2(n30070), .O(n27325) );
  MUX2S U19200 ( .A(n30044), .B(n30070), .S(gray_img[145]), .O(n27326) );
  AO12S U19201 ( .B1(n27821), .B2(n27820), .A1(n27819), .O(n13791) );
  ND2S U19202 ( .I1(n15929), .I2(n27814), .O(n27815) );
  MUX2S U19203 ( .A(n30005), .B(n27814), .S(gray_img[25]), .O(n27816) );
  AO12S U19204 ( .B1(n29904), .B2(n29893), .A1(n29892), .O(n13975) );
  ND2S U19205 ( .I1(n15929), .I2(n29898), .O(n29889) );
  MUX2S U19206 ( .A(n29566), .B(n29898), .S(gray_img[649]), .O(n29890) );
  AO12S U19207 ( .B1(n28950), .B2(n28949), .A1(n28948), .O(n14045) );
  ND2S U19208 ( .I1(n15932), .I2(n28943), .O(n28944) );
  MUX2S U19209 ( .A(n29032), .B(n28943), .S(gray_img[537]), .O(n28945) );
  OA12S U19210 ( .B1(n29884), .B2(n29883), .A1(n29882), .O(n29885) );
  MUX2S U19211 ( .A(n30005), .B(n29881), .S(gray_img[521]), .O(n29882) );
  AO12S U19212 ( .B1(n27840), .B2(n26296), .A1(n26295), .O(n14106) );
  ND2S U19213 ( .I1(n15885), .I2(n27834), .O(n26292) );
  MUX2S U19214 ( .A(n29566), .B(n27834), .S(gray_img[433]), .O(n26293) );
  OA12S U19215 ( .B1(n29884), .B2(n27224), .A1(n27223), .O(n27228) );
  ND2S U19216 ( .I1(n27226), .I2(n27225), .O(n27227) );
  MUX2S U19217 ( .A(n30056), .B(n27222), .S(gray_img[417]), .O(n27223) );
  OA12S U19218 ( .B1(n29884), .B2(n27254), .A1(n27253), .O(n27255) );
  ND2S U19219 ( .I1(n27251), .I2(n27250), .O(n27256) );
  MUX2S U19220 ( .A(n30050), .B(n27252), .S(gray_img[289]), .O(n27253) );
  AO12S U19221 ( .B1(n27785), .B2(n27517), .A1(n27516), .O(n14194) );
  ND2S U19222 ( .I1(n15931), .I2(n27779), .O(n27513) );
  MUX2S U19223 ( .A(n29597), .B(n27779), .S(gray_img[177]), .O(n27514) );
  AO12S U19224 ( .B1(n27708), .B2(n27697), .A1(n27696), .O(n14229) );
  MUX2S U19225 ( .A(n30005), .B(n27702), .S(gray_img[57]), .O(n27694) );
  AO12S U19226 ( .B1(n26931), .B2(n26930), .A1(n26929), .O(n14256) );
  ND2S U19227 ( .I1(n15931), .I2(n26924), .O(n26925) );
  MUX2S U19228 ( .A(n30056), .B(n26924), .S(gray_img[33]), .O(n26926) );
  AO12S U19229 ( .B1(n29350), .B2(n28919), .A1(n28918), .O(n14268) );
  ND2S U19230 ( .I1(n15931), .I2(n29344), .O(n28915) );
  MUX2S U19231 ( .A(n30005), .B(n29344), .S(gray_img[665]), .O(n28916) );
  AO12S U19232 ( .B1(n15885), .B2(n25473), .A1(n25472), .O(n14281) );
  AO12S U19233 ( .B1(n15884), .B2(n25761), .A1(n25461), .O(n14282) );
  AO12S U19234 ( .B1(n15885), .B2(n28803), .A1(n25632), .O(n14283) );
  ND2S U19235 ( .I1(n15931), .I2(n20202), .O(n18783) );
  ND2S U19236 ( .I1(n15931), .I2(n20586), .O(n20587) );
  ND2S U19237 ( .I1(n15931), .I2(n20424), .O(n18840) );
  MUX2S U19238 ( .A(n20842), .B(n20424), .S(gray_img[1929]), .O(n18839) );
  ND2S U19239 ( .I1(n15931), .I2(n20063), .O(n18503) );
  MUX2S U19240 ( .A(n29597), .B(n20063), .S(gray_img[1905]), .O(n18502) );
  ND2S U19241 ( .I1(n15931), .I2(n20544), .O(n20546) );
  MUX2S U19242 ( .A(n30050), .B(n20544), .S(gray_img[1897]), .O(n20545) );
  AO12S U19243 ( .B1(n15884), .B2(n25832), .A1(n25825), .O(n14296) );
  MUX2S U19244 ( .A(n27447), .B(n25830), .S(gray_img[1889]), .O(n25825) );
  AO12S U19245 ( .B1(n15884), .B2(n25477), .A1(n25474), .O(n14297) );
  MUX2S U19246 ( .A(n27447), .B(n25475), .S(gray_img[1881]), .O(n25474) );
  AO12S U19247 ( .B1(n15884), .B2(n25460), .A1(n25459), .O(n14298) );
  MUX2S U19248 ( .A(n27447), .B(n25458), .S(gray_img[1873]), .O(n25459) );
  AO12S U19249 ( .B1(n15884), .B2(n25631), .A1(n25630), .O(n14299) );
  MUX2S U19250 ( .A(n27447), .B(n25629), .S(gray_img[1865]), .O(n25630) );
  MUX2S U19251 ( .A(n29587), .B(n20142), .S(gray_img[1833]), .O(n19595) );
  ND2S U19252 ( .I1(n15931), .I2(n20319), .O(n18844) );
  MUX2S U19253 ( .A(n20808), .B(n20319), .S(gray_img[1801]), .O(n18843) );
  MUX2S U19254 ( .A(n30044), .B(n20449), .S(gray_img[1769]), .O(n19536) );
  AO12S U19255 ( .B1(n15884), .B2(n25510), .A1(n25509), .O(n14313) );
  AO12S U19256 ( .B1(n15885), .B2(n25498), .A1(n25495), .O(n14314) );
  MUX2S U19257 ( .A(n28534), .B(n25496), .S(gray_img[1745]), .O(n25495) );
  AO12S U19258 ( .B1(n15885), .B2(n25649), .A1(n25648), .O(n14315) );
  MUX2S U19259 ( .A(n15889), .B(n25647), .S(gray_img[1737]), .O(n25648) );
  MUX2S U19260 ( .A(n29566), .B(n19955), .S(gray_img[1729]), .O(n19528) );
  ND2S U19261 ( .I1(n15931), .I2(n20509), .O(n18796) );
  MUX2S U19262 ( .A(n25928), .B(n20509), .S(gray_img[1657]), .O(n18795) );
  ND2S U19263 ( .I1(n15885), .I2(n20525), .O(n18501) );
  MUX2S U19264 ( .A(n29587), .B(n20525), .S(gray_img[1649]), .O(n18500) );
  AO12S U19265 ( .B1(n15884), .B2(n25576), .A1(n25511), .O(n14329) );
  MUX2S U19266 ( .A(n27447), .B(n25574), .S(gray_img[1625]), .O(n25511) );
  AO12S U19267 ( .B1(n15928), .B2(n25494), .A1(n25487), .O(n14330) );
  ND2S U19268 ( .I1(n15885), .I2(n20731), .O(n20690) );
  MUX2S U19269 ( .A(n30050), .B(n20731), .S(gray_img[1593]), .O(n20689) );
  ND2S U19270 ( .I1(n15885), .I2(n20839), .O(n20771) );
  MUX2S U19271 ( .A(n20830), .B(n20839), .S(gray_img[1585]), .O(n20772) );
  ND2S U19272 ( .I1(n15885), .I2(n20395), .O(n19654) );
  MUX2S U19273 ( .A(n30050), .B(n20395), .S(gray_img[1577]), .O(n19655) );
  ND2S U19274 ( .I1(n15885), .I2(n20824), .O(n19652) );
  MUX2S U19275 ( .A(n30056), .B(n20824), .S(gray_img[1569]), .O(n19653) );
  MUX2S U19276 ( .A(n30044), .B(n20596), .S(gray_img[1561]), .O(n19543) );
  MUX2S U19277 ( .A(n29566), .B(n20602), .S(gray_img[1553]), .O(n19549) );
  MUX2S U19278 ( .A(n29587), .B(n20550), .S(gray_img[1545]), .O(n19516) );
  MUX2S U19279 ( .A(n20808), .B(n20512), .S(gray_img[1521]), .O(n19514) );
  AO12S U19280 ( .B1(n15932), .B2(n27971), .A1(n27970), .O(n14344) );
  AO12S U19281 ( .B1(n15884), .B2(n28355), .A1(n28354), .O(n14345) );
  ND2S U19282 ( .I1(n15885), .I2(n20821), .O(n20822) );
  MUX2S U19283 ( .A(n30044), .B(n20821), .S(gray_img[1457]), .O(n20823) );
  MUX2S U19284 ( .A(n30044), .B(n20293), .S(gray_img[1433]), .O(n19569) );
  MUX2S U19285 ( .A(n20842), .B(n20193), .S(gray_img[1425]), .O(n19571) );
  ND2S U19286 ( .I1(n15885), .I2(n20035), .O(n18722) );
  MUX2S U19287 ( .A(n20842), .B(n20035), .S(gray_img[1417]), .O(n18721) );
  MUX2S U19288 ( .A(n30056), .B(n20571), .S(gray_img[1401]), .O(n19502) );
  ND2S U19289 ( .I1(n15885), .I2(n20722), .O(n20724) );
  MUX2S U19290 ( .A(n30050), .B(n20722), .S(gray_img[1385]), .O(n20723) );
  AO12S U19291 ( .B1(n15885), .B2(n28203), .A1(n27972), .O(n14360) );
  MUX2S U19292 ( .A(n28534), .B(n28201), .S(gray_img[1377]), .O(n27972) );
  AO12S U19293 ( .B1(n15884), .B2(n28536), .A1(n28535), .O(n14363) );
  MUX2S U19294 ( .A(n28534), .B(n28533), .S(gray_img[1353]), .O(n28535) );
  ND2S U19295 ( .I1(n15885), .I2(n20734), .O(n20736) );
  MUX2S U19296 ( .A(n29597), .B(n20734), .S(gray_img[1345]), .O(n20735) );
  ND2S U19297 ( .I1(n15885), .I2(n20833), .O(n20834) );
  MUX2S U19298 ( .A(n30044), .B(n20833), .S(gray_img[1329]), .O(n20835) );
  MUX2S U19299 ( .A(n30056), .B(n20362), .S(gray_img[1297]), .O(n19593) );
  ND2S U19300 ( .I1(n15885), .I2(n20725), .O(n20727) );
  MUX2S U19301 ( .A(n20808), .B(n20725), .S(gray_img[1265]), .O(n20726) );
  AO12S U19302 ( .B1(n15931), .B2(n28288), .A1(n28285), .O(n14377) );
  AO12S U19303 ( .B1(n15885), .B2(n28271), .A1(n28270), .O(n14378) );
  AO12S U19304 ( .B1(n15884), .B2(n28475), .A1(n28474), .O(n14379) );
  AO12S U19305 ( .B1(n15885), .B2(n28092), .A1(n28023), .O(n14392) );
  AO12S U19306 ( .B1(n15884), .B2(n28284), .A1(n28277), .O(n14393) );
  AO12S U19307 ( .B1(n15884), .B2(n28480), .A1(n28476), .O(n14395) );
  ND2S U19308 ( .I1(n20752), .I2(n20751), .O(n14397) );
  ND2S U19309 ( .I1(n15885), .I2(n20760), .O(n20752) );
  MUX2S U19310 ( .A(n30056), .B(n20760), .S(gray_img[1081]), .O(n20751) );
  ND2S U19311 ( .I1(n15885), .I2(n20854), .O(n20852) );
  MUX2S U19312 ( .A(n30044), .B(n20854), .S(gray_img[1073]), .O(n20853) );
  ND2S U19313 ( .I1(n15885), .I2(n20368), .O(n18512) );
  MUX2S U19314 ( .A(n15904), .B(n20368), .S(gray_img[1057]), .O(n18513) );
  MUX2S U19315 ( .A(n15904), .B(n20562), .S(gray_img[1009]), .O(n19484) );
  ND2S U19316 ( .I1(n15885), .I2(n20384), .O(n18921) );
  ND2S U19317 ( .I1(n15885), .I2(n20580), .O(n20581) );
  MUX2S U19318 ( .A(n29587), .B(n20580), .S(gray_img[961]), .O(n20582) );
  MUX2S U19319 ( .A(n30005), .B(n20559), .S(gray_img[881]), .O(n19482) );
  ND2S U19320 ( .I1(n15885), .I2(n20212), .O(n18915) );
  MUX2S U19321 ( .A(n30005), .B(n20212), .S(gray_img[873]), .O(n18916) );
  AO12S U19322 ( .B1(n15933), .B2(n27190), .A1(n27189), .O(n14419) );
  ND2S U19323 ( .I1(n15885), .I2(n20365), .O(n18917) );
  MUX2S U19324 ( .A(n30005), .B(n20365), .S(gray_img[745]), .O(n18918) );
  AO12S U19325 ( .B1(n15884), .B2(n26155), .A1(n26154), .O(n14424) );
  MUX2S U19326 ( .A(n27447), .B(n26153), .S(gray_img[737]), .O(n26154) );
  AO12S U19327 ( .B1(n15884), .B2(n26160), .A1(n26156), .O(n14432) );
  AO12S U19328 ( .B1(n15885), .B2(n27133), .A1(n27132), .O(n14435) );
  MUX2S U19329 ( .A(n29597), .B(n20480), .S(gray_img[489]), .O(n19808) );
  MUX2S U19330 ( .A(n25928), .B(n20486), .S(gray_img[377]), .O(n19480) );
  AO12S U19331 ( .B1(n15884), .B2(n26861), .A1(n26860), .O(n14451) );
  MUX2S U19332 ( .A(n15889), .B(n26859), .S(gray_img[329]), .O(n26860) );
  ND2S U19333 ( .I1(n15885), .I2(n20620), .O(n20622) );
  MUX2S U19334 ( .A(n30044), .B(n20620), .S(gray_img[233]), .O(n20621) );
  AO12S U19335 ( .B1(n15886), .B2(n26883), .A1(n26880), .O(n14459) );
  ND2S U19336 ( .I1(n15884), .I2(n20617), .O(n20619) );
  MUX2S U19337 ( .A(n29587), .B(n20617), .S(gray_img[105]), .O(n20618) );
  ND2S U19338 ( .I1(n22655), .I2(n22654), .O(n15814) );
  AO12S U19339 ( .B1(n28847), .B2(n28800), .A1(n28799), .O(n14475) );
  ND2S U19340 ( .I1(n15937), .I2(n28840), .O(n28796) );
  MUX2S U19341 ( .A(n15904), .B(n28840), .S(gray_img[138]), .O(n28797) );
  ND2S U19342 ( .I1(n28727), .I2(n28231), .O(n28234) );
  OA12S U19343 ( .B1(n29849), .B2(n28730), .A1(n28232), .O(n28233) );
  MUX2S U19344 ( .A(n15904), .B(n28728), .S(gray_img[410]), .O(n28232) );
  AO12S U19345 ( .B1(n28724), .B2(n26072), .A1(n26071), .O(n13656) );
  ND2S U19346 ( .I1(n15883), .I2(n28718), .O(n26068) );
  MUX2S U19347 ( .A(n15904), .B(n28718), .S(gray_img[954]), .O(n26069) );
  AO12S U19348 ( .B1(n26096), .B2(n25927), .A1(n25926), .O(n13657) );
  ND2S U19349 ( .I1(n15934), .I2(n26090), .O(n25923) );
  MUX2S U19350 ( .A(n15904), .B(n26090), .S(gray_img[946]), .O(n25924) );
  ND2S U19351 ( .I1(n28806), .I2(n28700), .O(n28703) );
  MUX2S U19352 ( .A(n29587), .B(n28807), .S(gray_img[402]), .O(n28701) );
  AO12S U19353 ( .B1(n25619), .B2(n25602), .A1(n25601), .O(n13658) );
  ND2S U19354 ( .I1(n15934), .I2(n25612), .O(n25598) );
  MUX2S U19355 ( .A(n30056), .B(n25612), .S(gray_img[938]), .O(n25599) );
  AO12S U19356 ( .B1(n25758), .B2(n25739), .A1(n25738), .O(n13659) );
  ND2S U19357 ( .I1(n15935), .I2(n25751), .O(n25735) );
  MUX2S U19358 ( .A(n30050), .B(n25751), .S(gray_img[930]), .O(n25736) );
  AO12S U19359 ( .B1(n30128), .B2(n30062), .A1(n30061), .O(n14476) );
  ND2S U19360 ( .I1(n15937), .I2(n30121), .O(n30058) );
  MUX2S U19361 ( .A(n30056), .B(n30121), .S(gray_img[130]), .O(n30059) );
  AO12S U19362 ( .B1(n30038), .B2(n29373), .A1(n29372), .O(n14473) );
  ND2S U19363 ( .I1(n15935), .I2(n30032), .O(n29369) );
  MUX2S U19364 ( .A(n30044), .B(n30032), .S(gray_img[394]), .O(n29370) );
  MUX2S U19365 ( .A(n30044), .B(n23195), .S(gray_img[922]), .O(n23174) );
  ND2S U19366 ( .I1(n30020), .I2(n29177), .O(n29180) );
  OA12S U19367 ( .B1(n29849), .B2(n30023), .A1(n29178), .O(n29179) );
  MUX2S U19368 ( .A(n15904), .B(n30021), .S(gray_img[914]), .O(n29178) );
  AO12S U19369 ( .B1(n30109), .B2(n29990), .A1(n29989), .O(n14474) );
  ND2S U19370 ( .I1(n15937), .I2(n30103), .O(n29986) );
  MUX2S U19371 ( .A(n30050), .B(n30103), .S(gray_img[386]), .O(n29987) );
  AO12S U19372 ( .B1(n29604), .B2(n29576), .A1(n29575), .O(n13662) );
  ND2S U19373 ( .I1(n15936), .I2(n29598), .O(n29572) );
  MUX2S U19374 ( .A(n29597), .B(n29598), .S(gray_img[906]), .O(n29573) );
  AO12S U19375 ( .B1(n30098), .B2(n29476), .A1(n29475), .O(n13663) );
  ND2S U19376 ( .I1(n15937), .I2(n30092), .O(n29472) );
  MUX2S U19377 ( .A(n29597), .B(n30092), .S(gray_img[898]), .O(n29473) );
  AO12S U19378 ( .B1(n26080), .B2(n26044), .A1(n26043), .O(n13664) );
  ND2S U19379 ( .I1(n15937), .I2(n26073), .O(n26040) );
  MUX2S U19380 ( .A(n15904), .B(n26073), .S(gray_img[826]), .O(n26041) );
  AO12S U19381 ( .B1(n25936), .B2(n25896), .A1(n25895), .O(n13665) );
  MUX2S U19382 ( .A(n25928), .B(n25929), .S(gray_img[818]), .O(n25893) );
  OA12S U19383 ( .B1(n29849), .B2(n25607), .A1(n25570), .O(n25571) );
  MUX2S U19384 ( .A(n25928), .B(n25605), .S(gray_img[810]), .O(n25570) );
  AO12S U19385 ( .B1(n25750), .B2(n25714), .A1(n25713), .O(n13667) );
  ND2S U19386 ( .I1(n15937), .I2(n25744), .O(n25710) );
  MUX2S U19387 ( .A(n25928), .B(n25744), .S(gray_img[802]), .O(n25711) );
  AO12S U19388 ( .B1(n29273), .B2(n29257), .A1(n29256), .O(n13668) );
  ND2S U19389 ( .I1(n15937), .I2(n29266), .O(n29253) );
  MUX2S U19390 ( .A(n30056), .B(n29266), .S(gray_img[794]), .O(n29254) );
  AO12S U19391 ( .B1(n29192), .B2(n29156), .A1(n29155), .O(n13669) );
  ND2S U19392 ( .I1(n15937), .I2(n29186), .O(n29152) );
  MUX2S U19393 ( .A(n30056), .B(n29186), .S(gray_img[786]), .O(n29153) );
  AO12S U19394 ( .B1(n29487), .B2(n29451), .A1(n29450), .O(n13671) );
  MUX2S U19395 ( .A(n30050), .B(n29481), .S(gray_img[770]), .O(n29448) );
  ND2S U19396 ( .I1(n28247), .I2(n28196), .O(n28199) );
  OA12S U19397 ( .B1(n29849), .B2(n28250), .A1(n28197), .O(n28198) );
  MUX2S U19398 ( .A(n30005), .B(n28248), .S(gray_img[282]), .O(n28197) );
  ND2S U19399 ( .I1(n28136), .I2(n27949), .O(n27952) );
  OA12S U19400 ( .B1(n29849), .B2(n28139), .A1(n27950), .O(n27951) );
  MUX2S U19401 ( .A(n30005), .B(n28137), .S(gray_img[698]), .O(n27950) );
  AO12S U19402 ( .B1(n28214), .B2(n28120), .A1(n28119), .O(n13673) );
  ND2S U19403 ( .I1(n15937), .I2(n28208), .O(n28116) );
  MUX2S U19404 ( .A(n30005), .B(n28208), .S(gray_img[690]), .O(n28117) );
  OA12S U19405 ( .B1(n29849), .B2(n28709), .A1(n28665), .O(n28666) );
  MUX2S U19406 ( .A(n30050), .B(n28707), .S(gray_img[274]), .O(n28665) );
  AO12S U19407 ( .B1(n29381), .B2(n29339), .A1(n29338), .O(n13705) );
  ND2S U19408 ( .I1(n15934), .I2(n29374), .O(n29335) );
  MUX2S U19409 ( .A(n29597), .B(n29374), .S(gray_img[266]), .O(n29336) );
  AO12S U19410 ( .B1(n30012), .B2(n29965), .A1(n29964), .O(n13734) );
  ND2S U19411 ( .I1(n15936), .I2(n30006), .O(n29961) );
  MUX2S U19412 ( .A(n15904), .B(n30006), .S(gray_img[258]), .O(n29962) );
  AO12S U19413 ( .B1(n30087), .B2(n28839), .A1(n28838), .O(n13752) );
  ND2S U19414 ( .I1(n15937), .I2(n30081), .O(n28835) );
  MUX2S U19415 ( .A(n30044), .B(n30081), .S(gray_img[10]), .O(n28836) );
  AO12S U19416 ( .B1(n27851), .B2(n27813), .A1(n27812), .O(n13760) );
  ND2S U19417 ( .I1(n15937), .I2(n27845), .O(n27809) );
  MUX2S U19418 ( .A(n29587), .B(n27845), .S(gray_img[154]), .O(n27810) );
  AO12S U19419 ( .B1(n30076), .B2(n27324), .A1(n27323), .O(n13770) );
  ND2S U19420 ( .I1(n15937), .I2(n30070), .O(n27320) );
  MUX2S U19421 ( .A(n30044), .B(n30070), .S(gray_img[146]), .O(n27321) );
  AO12S U19422 ( .B1(n27821), .B2(n27771), .A1(n27770), .O(n13790) );
  ND2S U19423 ( .I1(n15934), .I2(n27814), .O(n27767) );
  MUX2S U19424 ( .A(n30005), .B(n27814), .S(gray_img[26]), .O(n27768) );
  AO12S U19425 ( .B1(n27378), .B2(n27349), .A1(n27348), .O(n13800) );
  ND2S U19426 ( .I1(n15934), .I2(n27371), .O(n27345) );
  MUX2S U19427 ( .A(n30005), .B(n27371), .S(gray_img[18]), .O(n27346) );
  AO12S U19428 ( .B1(n28588), .B2(n28557), .A1(n28556), .O(n13949) );
  ND2S U19429 ( .I1(n15934), .I2(n28581), .O(n28553) );
  MUX2S U19430 ( .A(n30050), .B(n28581), .S(gray_img[674]), .O(n28554) );
  AO12S U19431 ( .B1(n29350), .B2(n28914), .A1(n28913), .O(n13957) );
  ND2S U19432 ( .I1(n15883), .I2(n29344), .O(n28910) );
  MUX2S U19433 ( .A(n30056), .B(n29344), .S(gray_img[666]), .O(n28911) );
  AO12S U19434 ( .B1(n29040), .B2(n29008), .A1(n29007), .O(n13965) );
  ND2S U19435 ( .I1(n15937), .I2(n29033), .O(n29004) );
  MUX2S U19436 ( .A(n29597), .B(n29033), .S(gray_img[658]), .O(n29005) );
  AO12S U19437 ( .B1(n29904), .B2(n29878), .A1(n29877), .O(n13974) );
  ND2S U19438 ( .I1(n15935), .I2(n29898), .O(n29874) );
  MUX2S U19439 ( .A(n30050), .B(n29898), .S(gray_img[650]), .O(n29875) );
  ND2S U19440 ( .I1(n29993), .I2(n29701), .O(n29704) );
  OA12S U19441 ( .B1(n29849), .B2(n29996), .A1(n29702), .O(n29703) );
  MUX2S U19442 ( .A(n15904), .B(n29994), .S(gray_img[642]), .O(n29702) );
  ND2S U19443 ( .I1(n23492), .I2(n23335), .O(n23338) );
  MUX2S U19444 ( .A(n30050), .B(n23493), .S(gray_img[570]), .O(n23336) );
  AO12S U19445 ( .B1(n28128), .B2(n28089), .A1(n28088), .O(n14017) );
  ND2S U19446 ( .I1(n15937), .I2(n28121), .O(n28085) );
  MUX2S U19447 ( .A(n30044), .B(n28121), .S(gray_img[562]), .O(n28086) );
  AO12S U19448 ( .B1(n28459), .B2(n28420), .A1(n28419), .O(n14026) );
  ND2S U19449 ( .I1(n15934), .I2(n28452), .O(n28416) );
  MUX2S U19450 ( .A(n29032), .B(n28452), .S(gray_img[554]), .O(n28417) );
  ND2S U19451 ( .I1(n28671), .I2(n28576), .O(n28579) );
  OA12S U19452 ( .B1(n29849), .B2(n28674), .A1(n28577), .O(n28578) );
  MUX2S U19453 ( .A(n15904), .B(n28672), .S(gray_img[546]), .O(n28577) );
  AO12S U19454 ( .B1(n28950), .B2(n28934), .A1(n28933), .O(n14044) );
  ND2S U19455 ( .I1(n15937), .I2(n28943), .O(n28930) );
  MUX2S U19456 ( .A(n29032), .B(n28943), .S(gray_img[538]), .O(n28931) );
  OA12S U19457 ( .B1(n29849), .B2(n29883), .A1(n29848), .O(n29850) );
  MUX2S U19458 ( .A(n30005), .B(n29881), .S(gray_img[522]), .O(n29848) );
  OA12S U19459 ( .B1(n29849), .B2(n29742), .A1(n29727), .O(n29728) );
  MUX2S U19460 ( .A(n15904), .B(n29740), .S(gray_img[514]), .O(n29727) );
  AO12S U19461 ( .B1(n26473), .B2(n26436), .A1(n26435), .O(n14096) );
  ND2S U19462 ( .I1(n15935), .I2(n26466), .O(n26432) );
  MUX2S U19463 ( .A(n30044), .B(n26466), .S(gray_img[442]), .O(n26433) );
  AO12S U19464 ( .B1(n27840), .B2(n26291), .A1(n26290), .O(n14105) );
  ND2S U19465 ( .I1(n15937), .I2(n27834), .O(n26287) );
  MUX2S U19466 ( .A(n15904), .B(n27834), .S(gray_img[434]), .O(n26288) );
  ND2S U19467 ( .I1(n23121), .I2(n23095), .O(n23098) );
  MUX2S U19468 ( .A(n29587), .B(n25151), .S(gray_img[426]), .O(n23096) );
  OA12S U19469 ( .B1(n29849), .B2(n27224), .A1(n27217), .O(n27220) );
  ND2S U19470 ( .I1(n27226), .I2(n27218), .O(n27219) );
  MUX2S U19471 ( .A(n30050), .B(n27222), .S(gray_img[418]), .O(n27217) );
  AO12S U19472 ( .B1(n26489), .B2(n26465), .A1(n26464), .O(n14140) );
  ND2S U19473 ( .I1(n15936), .I2(n26483), .O(n26461) );
  MUX2S U19474 ( .A(n15904), .B(n26483), .S(gray_img[314]), .O(n26462) );
  ND2S U19475 ( .I1(n26327), .I2(n26313), .O(n26314) );
  OA12S U19476 ( .B1(n29849), .B2(n26324), .A1(n26312), .O(n26315) );
  MUX2S U19477 ( .A(n15904), .B(n26322), .S(gray_img[306]), .O(n26312) );
  AO12S U19478 ( .B1(n27121), .B2(n27102), .A1(n27101), .O(n14158) );
  ND2S U19479 ( .I1(n15937), .I2(n27114), .O(n27098) );
  MUX2S U19480 ( .A(n29587), .B(n27114), .S(gray_img[298]), .O(n27099) );
  OA12S U19481 ( .B1(n29849), .B2(n27254), .A1(n27237), .O(n27238) );
  ND2S U19482 ( .I1(n27251), .I2(n27236), .O(n27239) );
  MUX2S U19483 ( .A(n29587), .B(n27252), .S(gray_img[290]), .O(n27237) );
  AO12S U19484 ( .B1(n27692), .B2(n27656), .A1(n27655), .O(n14184) );
  ND2S U19485 ( .I1(n15936), .I2(n27685), .O(n27652) );
  MUX2S U19486 ( .A(n30044), .B(n27685), .S(gray_img[186]), .O(n27653) );
  AO12S U19487 ( .B1(n27785), .B2(n27511), .A1(n27510), .O(n14193) );
  ND2S U19488 ( .I1(n15935), .I2(n27779), .O(n27507) );
  MUX2S U19489 ( .A(n30050), .B(n27779), .S(gray_img[178]), .O(n27508) );
  OA12S U19490 ( .B1(n29849), .B2(n27358), .A1(n26819), .O(n26820) );
  MUX2S U19491 ( .A(n30050), .B(n27356), .S(gray_img[170]), .O(n26819) );
  AO12S U19492 ( .B1(n26939), .B2(n26923), .A1(n26922), .O(n14211) );
  ND2S U19493 ( .I1(n15935), .I2(n26932), .O(n26919) );
  MUX2S U19494 ( .A(n29032), .B(n26932), .S(gray_img[162]), .O(n26920) );
  AO12S U19495 ( .B1(n27708), .B2(n27684), .A1(n27683), .O(n14228) );
  ND2S U19496 ( .I1(n15935), .I2(n27702), .O(n27680) );
  MUX2S U19497 ( .A(n30050), .B(n27702), .S(gray_img[58]), .O(n27681) );
  AO12S U19498 ( .B1(n27556), .B2(n27537), .A1(n27536), .O(n14237) );
  ND2S U19499 ( .I1(n15934), .I2(n27550), .O(n27533) );
  MUX2S U19500 ( .A(n29032), .B(n27550), .S(gray_img[50]), .O(n27534) );
  AO12S U19501 ( .B1(n26849), .B2(n26838), .A1(n26837), .O(n14246) );
  ND2S U19502 ( .I1(n15935), .I2(n26842), .O(n26834) );
  MUX2S U19503 ( .A(n30050), .B(n26842), .S(gray_img[42]), .O(n26835) );
  AO12S U19504 ( .B1(n26931), .B2(n26903), .A1(n26902), .O(n14255) );
  ND2S U19505 ( .I1(n15937), .I2(n26924), .O(n26899) );
  MUX2S U19506 ( .A(n29587), .B(n26924), .S(gray_img[34]), .O(n26900) );
  AO12S U19507 ( .B1(n28607), .B2(n28451), .A1(n28450), .O(n14470) );
  ND2S U19508 ( .I1(n15935), .I2(n28601), .O(n28447) );
  MUX2S U19509 ( .A(n15904), .B(n28601), .S(gray_img[682]), .O(n28448) );
  AO12S U19510 ( .B1(n15883), .B2(n25836), .A1(n25829), .O(n14481) );
  AO12S U19511 ( .B1(n15882), .B2(n25473), .A1(n25465), .O(n14482) );
  AO12S U19512 ( .B1(n15883), .B2(n25761), .A1(n25457), .O(n14483) );
  AO12S U19513 ( .B1(n15883), .B2(n28803), .A1(n25628), .O(n14484) );
  ND2S U19514 ( .I1(n15937), .I2(n20209), .O(n18945) );
  ND2S U19515 ( .I1(n15937), .I2(n20849), .O(n20792) );
  MUX2S U19516 ( .A(n29597), .B(n20849), .S(gray_img[1970]), .O(n20793) );
  MUX2S U19517 ( .A(n29587), .B(n19970), .S(gray_img[1946]), .O(n19615) );
  MUX2S U19518 ( .A(n29587), .B(n20389), .S(gray_img[1938]), .O(n19627) );
  MUX2S U19519 ( .A(n20808), .B(n20424), .S(gray_img[1930]), .O(n19476) );
  MUX2S U19520 ( .A(n30050), .B(n20430), .S(gray_img[1914]), .O(n19474) );
  MUX2S U19521 ( .A(n30056), .B(n20544), .S(gray_img[1898]), .O(n19470) );
  AO12S U19522 ( .B1(n15938), .B2(n25832), .A1(n25824), .O(n14497) );
  AO12S U19523 ( .B1(n15934), .B2(n25477), .A1(n25470), .O(n14498) );
  AO12S U19524 ( .B1(n15938), .B2(n25460), .A1(n25453), .O(n14499) );
  MUX2S U19525 ( .A(n28534), .B(n25458), .S(gray_img[1874]), .O(n25453) );
  AO12S U19526 ( .B1(n15938), .B2(n25631), .A1(n25623), .O(n14500) );
  MUX2S U19527 ( .A(n15889), .B(n25629), .S(gray_img[1866]), .O(n25623) );
  MUX2S U19528 ( .A(n29597), .B(n20504), .S(gray_img[1858]), .O(n19468) );
  ND2S U19529 ( .I1(n15937), .I2(n20740), .O(n20671) );
  MUX2S U19530 ( .A(n29597), .B(n20740), .S(gray_img[1850]), .O(n20670) );
  ND2S U19531 ( .I1(n15937), .I2(n20862), .O(n20863) );
  MUX2S U19532 ( .A(n29597), .B(n20862), .S(gray_img[1842]), .O(n20864) );
  ND2S U19533 ( .I1(n15937), .I2(n20142), .O(n18781) );
  MUX2S U19534 ( .A(n29566), .B(n20142), .S(gray_img[1834]), .O(n18782) );
  MUX2S U19535 ( .A(n29587), .B(n20296), .S(gray_img[1818]), .O(n19591) );
  MUX2S U19536 ( .A(n29566), .B(n20354), .S(gray_img[1810]), .O(n20343) );
  MUX2S U19537 ( .A(n20842), .B(n20319), .S(gray_img[1802]), .O(n19460) );
  ND2S U19538 ( .I1(n15937), .I2(n20547), .O(n20549) );
  MUX2S U19539 ( .A(n29597), .B(n20547), .S(gray_img[1786]), .O(n20548) );
  ND2S U19540 ( .I1(n15937), .I2(n20541), .O(n20543) );
  MUX2S U19541 ( .A(n29597), .B(n20541), .S(gray_img[1778]), .O(n20542) );
  MUX2S U19542 ( .A(n30050), .B(n20449), .S(gray_img[1770]), .O(n19458) );
  AO12S U19543 ( .B1(n15939), .B2(n25778), .A1(n25770), .O(n14513) );
  MUX2S U19544 ( .A(n27447), .B(n25776), .S(gray_img[1762]), .O(n25770) );
  AO12S U19545 ( .B1(n15883), .B2(n25510), .A1(n25502), .O(n14514) );
  MUX2S U19546 ( .A(n15889), .B(n25508), .S(gray_img[1754]), .O(n25502) );
  AO12S U19547 ( .B1(n15883), .B2(n25498), .A1(n25491), .O(n14515) );
  AO12S U19548 ( .B1(n15883), .B2(n25649), .A1(n25641), .O(n14516) );
  MUX2S U19549 ( .A(n15889), .B(n25647), .S(gray_img[1738]), .O(n25641) );
  MUX2S U19550 ( .A(n29597), .B(n19955), .S(gray_img[1730]), .O(n19454) );
  ND2S U19551 ( .I1(n15937), .I2(n20737), .O(n20739) );
  MUX2S U19552 ( .A(n30044), .B(n20737), .S(gray_img[1722]), .O(n20738) );
  ND2S U19553 ( .I1(n15938), .I2(n20846), .O(n20831) );
  MUX2S U19554 ( .A(n20830), .B(n20846), .S(gray_img[1714]), .O(n20832) );
  ND2S U19555 ( .I1(n15882), .I2(n20827), .O(n20828) );
  MUX2S U19556 ( .A(n30050), .B(n20827), .S(gray_img[1706]), .O(n20829) );
  ND2S U19557 ( .I1(n15882), .I2(n20787), .O(n19658) );
  MUX2S U19558 ( .A(n30056), .B(n20787), .S(gray_img[1698]), .O(n19659) );
  ND2S U19559 ( .I1(n15882), .I2(n20599), .O(n20589) );
  ND2S U19560 ( .I1(n15938), .I2(n20605), .O(n20578) );
  MUX2S U19561 ( .A(n30056), .B(n20605), .S(gray_img[1682]), .O(n20579) );
  ND2S U19562 ( .I1(n15938), .I2(n20531), .O(n20533) );
  MUX2S U19563 ( .A(n29566), .B(n20531), .S(gray_img[1674]), .O(n20532) );
  ND2S U19564 ( .I1(n15882), .I2(n20583), .O(n20584) );
  MUX2S U19565 ( .A(n29587), .B(n20583), .S(gray_img[1666]), .O(n20585) );
  ND2S U19566 ( .I1(n15934), .I2(n20509), .O(n20511) );
  MUX2S U19567 ( .A(n29587), .B(n20509), .S(gray_img[1658]), .O(n20510) );
  ND2S U19568 ( .I1(n15934), .I2(n20525), .O(n20527) );
  MUX2S U19569 ( .A(n29587), .B(n20525), .S(gray_img[1650]), .O(n20526) );
  MUX2S U19570 ( .A(n29587), .B(n20463), .S(gray_img[1642]), .O(n19452) );
  AO12S U19571 ( .B1(n15883), .B2(n25899), .A1(n25775), .O(n14529) );
  MUX2S U19572 ( .A(n27447), .B(n25897), .S(gray_img[1634]), .O(n25775) );
  AO12S U19573 ( .B1(n15938), .B2(n25576), .A1(n25507), .O(n14530) );
  AO12S U19574 ( .B1(n15882), .B2(n25494), .A1(n25486), .O(n14531) );
  AO12S U19575 ( .B1(n15937), .B2(n25653), .A1(n25646), .O(n14532) );
  MUX2S U19576 ( .A(n25928), .B(n20528), .S(gray_img[1602]), .O(n19448) );
  ND2S U19577 ( .I1(n15937), .I2(n20731), .O(n20665) );
  MUX2S U19578 ( .A(n30056), .B(n20731), .S(gray_img[1594]), .O(n20664) );
  ND2S U19579 ( .I1(n15882), .I2(n20839), .O(n20802) );
  MUX2S U19580 ( .A(n20830), .B(n20839), .S(gray_img[1586]), .O(n20803) );
  ND2S U19581 ( .I1(n15882), .I2(n20395), .O(n19660) );
  MUX2S U19582 ( .A(n30050), .B(n20395), .S(gray_img[1578]), .O(n19661) );
  ND2S U19583 ( .I1(n15882), .I2(n20824), .O(n20796) );
  MUX2S U19584 ( .A(n30056), .B(n20824), .S(gray_img[1570]), .O(n20797) );
  ND2S U19585 ( .I1(n15882), .I2(n20596), .O(n20574) );
  MUX2S U19586 ( .A(n29587), .B(n20596), .S(gray_img[1562]), .O(n20575) );
  ND2S U19587 ( .I1(n15882), .I2(n20602), .O(n20603) );
  MUX2S U19588 ( .A(n29566), .B(n20602), .S(gray_img[1554]), .O(n20604) );
  ND2S U19589 ( .I1(n15882), .I2(n20550), .O(n20521) );
  MUX2S U19590 ( .A(n29566), .B(n20550), .S(gray_img[1546]), .O(n20520) );
  ND2S U19591 ( .I1(n15882), .I2(n20881), .O(n20869) );
  MUX2S U19592 ( .A(n29566), .B(n20881), .S(gray_img[1538]), .O(n20870) );
  MUX2S U19593 ( .A(n30044), .B(n20556), .S(gray_img[1530]), .O(n19446) );
  ND2S U19594 ( .I1(n15882), .I2(n20440), .O(n19639) );
  MUX2S U19595 ( .A(n30056), .B(n20440), .S(gray_img[1514]), .O(n19638) );
  AO12S U19596 ( .B1(n15883), .B2(n27971), .A1(n27964), .O(n14545) );
  AO12S U19597 ( .B1(n15939), .B2(n28355), .A1(n28347), .O(n14546) );
  MUX2S U19598 ( .A(n28534), .B(n28353), .S(gray_img[1498]), .O(n28347) );
  AO12S U19599 ( .B1(n15883), .B2(n28342), .A1(n28334), .O(n14547) );
  MUX2S U19600 ( .A(n27447), .B(n28340), .S(gray_img[1490]), .O(n28334) );
  AO12S U19601 ( .B1(n15937), .B2(n28560), .A1(n28532), .O(n14548) );
  MUX2S U19602 ( .A(n27447), .B(n28558), .S(gray_img[1482]), .O(n28532) );
  ND2S U19603 ( .I1(n15882), .I2(n20684), .O(n20650) );
  MUX2S U19604 ( .A(n29566), .B(n20684), .S(gray_img[1474]), .O(n20649) );
  ND2S U19605 ( .I1(n15882), .I2(n20709), .O(n20711) );
  ND2S U19606 ( .I1(n15938), .I2(n20821), .O(n20773) );
  MUX2S U19607 ( .A(n30044), .B(n20821), .S(gray_img[1458]), .O(n20774) );
  ND2S U19608 ( .I1(n15938), .I2(n20814), .O(n20777) );
  MUX2S U19609 ( .A(n29566), .B(n20814), .S(gray_img[1450]), .O(n20778) );
  ND2S U19610 ( .I1(n15938), .I2(n20811), .O(n20779) );
  ND2S U19611 ( .I1(n15938), .I2(n20293), .O(n18631) );
  MUX2S U19612 ( .A(n30050), .B(n20293), .S(gray_img[1434]), .O(n18632) );
  MUX2S U19613 ( .A(n20842), .B(n20193), .S(gray_img[1426]), .O(n19567) );
  ND2S U19614 ( .I1(n15938), .I2(n20035), .O(n18724) );
  MUX2S U19615 ( .A(n20842), .B(n20035), .S(gray_img[1418]), .O(n18723) );
  ND2S U19616 ( .I1(n15938), .I2(n20359), .O(n18864) );
  MUX2S U19617 ( .A(n20808), .B(n20359), .S(gray_img[1410]), .O(n18865) );
  MUX2S U19618 ( .A(n30050), .B(n20571), .S(gray_img[1402]), .O(n19440) );
  ND2S U19619 ( .I1(n15938), .I2(n20722), .O(n20659) );
  MUX2S U19620 ( .A(n30044), .B(n20722), .S(gray_img[1386]), .O(n20658) );
  AO12S U19621 ( .B1(n15939), .B2(n28203), .A1(n27968), .O(n14561) );
  MUX2S U19622 ( .A(n28534), .B(n28201), .S(gray_img[1378]), .O(n27968) );
  AO12S U19623 ( .B1(n15882), .B2(n28359), .A1(n28352), .O(n14562) );
  AO12S U19624 ( .B1(n15938), .B2(n28596), .A1(n28339), .O(n14563) );
  AO12S U19625 ( .B1(n15883), .B2(n28536), .A1(n28526), .O(n14564) );
  MUX2S U19626 ( .A(n28534), .B(n28533), .S(gray_img[1354]), .O(n28526) );
  ND2S U19627 ( .I1(n15938), .I2(n20734), .O(n20644) );
  MUX2S U19628 ( .A(n29587), .B(n20734), .S(gray_img[1346]), .O(n20643) );
  ND2S U19629 ( .I1(n15938), .I2(n20695), .O(n20683) );
  MUX2S U19630 ( .A(n30056), .B(n20695), .S(gray_img[1338]), .O(n20682) );
  ND2S U19631 ( .I1(n15938), .I2(n20833), .O(n20783) );
  MUX2S U19632 ( .A(n30050), .B(n20833), .S(gray_img[1330]), .O(n20784) );
  ND2S U19633 ( .I1(n15882), .I2(n20836), .O(n20790) );
  MUX2S U19634 ( .A(n29566), .B(n20836), .S(gray_img[1322]), .O(n20791) );
  ND2S U19635 ( .I1(n15882), .I2(n20843), .O(n20798) );
  MUX2S U19636 ( .A(n30044), .B(n20843), .S(gray_img[1314]), .O(n20799) );
  MUX2S U19637 ( .A(n30044), .B(n20362), .S(gray_img[1298]), .O(n19581) );
  ND2S U19638 ( .I1(n15882), .I2(n20427), .O(n18730) );
  ND2S U19639 ( .I1(n15882), .I2(n20392), .O(n18870) );
  MUX2S U19640 ( .A(n29597), .B(n20392), .S(gray_img[1282]), .O(n18871) );
  ND2S U19641 ( .I1(n15882), .I2(n20655), .O(n20654) );
  MUX2S U19642 ( .A(n20808), .B(n20655), .S(gray_img[1274]), .O(n20653) );
  ND2S U19643 ( .I1(n15882), .I2(n20725), .O(n20661) );
  MUX2S U19644 ( .A(n20808), .B(n20725), .S(gray_img[1266]), .O(n20660) );
  ND2S U19645 ( .I1(n15882), .I2(n20719), .O(n20663) );
  MUX2S U19646 ( .A(n30044), .B(n20719), .S(gray_img[1258]), .O(n20662) );
  AO12S U19647 ( .B1(n15939), .B2(n28031), .A1(n28027), .O(n14577) );
  AO12S U19648 ( .B1(n15883), .B2(n28288), .A1(n28281), .O(n14578) );
  AO12S U19649 ( .B1(n15882), .B2(n28271), .A1(n28263), .O(n14579) );
  AO12S U19650 ( .B1(n15882), .B2(n28475), .A1(n28469), .O(n14580) );
  ND2S U19651 ( .I1(n15882), .I2(n20702), .O(n20694) );
  MUX2S U19652 ( .A(n29566), .B(n20702), .S(gray_img[1218]), .O(n20693) );
  ND2S U19653 ( .I1(n20759), .I2(n20758), .O(n14582) );
  ND2S U19654 ( .I1(n15882), .I2(n20757), .O(n20759) );
  MUX2S U19655 ( .A(n30044), .B(n20757), .S(gray_img[1210]), .O(n20758) );
  ND2S U19656 ( .I1(n15882), .I2(n20857), .O(n20819) );
  MUX2S U19657 ( .A(n30044), .B(n20857), .S(gray_img[1202]), .O(n20820) );
  ND2S U19658 ( .I1(n15883), .I2(n20435), .O(n19685) );
  MUX2S U19659 ( .A(n29597), .B(n20435), .S(gray_img[1194]), .O(n19684) );
  MUX2S U19660 ( .A(n29597), .B(n20379), .S(gray_img[1186]), .O(n19553) );
  MUX2S U19661 ( .A(n29566), .B(n20553), .S(gray_img[1162]), .O(n19426) );
  MUX2S U19662 ( .A(n29566), .B(n20240), .S(gray_img[1154]), .O(n19700) );
  ND2S U19663 ( .I1(n15883), .I2(n20716), .O(n20718) );
  MUX2S U19664 ( .A(n30044), .B(n20716), .S(gray_img[1146]), .O(n20717) );
  ND2S U19665 ( .I1(n15883), .I2(n20124), .O(n19641) );
  MUX2S U19666 ( .A(n20808), .B(n20124), .S(gray_img[1138]), .O(n19640) );
  ND2S U19667 ( .I1(n15883), .I2(n20728), .O(n20730) );
  AO12S U19668 ( .B1(n15883), .B2(n28092), .A1(n28022), .O(n14593) );
  MUX2S U19669 ( .A(n27447), .B(n28090), .S(gray_img[1122]), .O(n28022) );
  AO12S U19670 ( .B1(n15939), .B2(n28284), .A1(n28276), .O(n14594) );
  AO12S U19671 ( .B1(n15883), .B2(n28423), .A1(n28268), .O(n14595) );
  AO12S U19672 ( .B1(n15938), .B2(n28480), .A1(n28472), .O(n14596) );
  ND2S U19673 ( .I1(n15883), .I2(n20743), .O(n20745) );
  MUX2S U19674 ( .A(n30050), .B(n20743), .S(gray_img[1090]), .O(n20744) );
  ND2S U19675 ( .I1(n20756), .I2(n20755), .O(n14598) );
  ND2S U19676 ( .I1(n15883), .I2(n20760), .O(n20756) );
  MUX2S U19677 ( .A(n30056), .B(n20760), .S(gray_img[1082]), .O(n20755) );
  ND2S U19678 ( .I1(n15883), .I2(n20854), .O(n20855) );
  MUX2S U19679 ( .A(n30044), .B(n20854), .S(gray_img[1074]), .O(n20856) );
  ND2S U19680 ( .I1(n15883), .I2(n20611), .O(n20613) );
  MUX2S U19681 ( .A(n29566), .B(n20611), .S(gray_img[1066]), .O(n20612) );
  MUX2S U19682 ( .A(n29566), .B(n20184), .S(gray_img[1050]), .O(n19603) );
  ND2S U19683 ( .I1(n19783), .I2(n19782), .O(n14603) );
  ND2S U19684 ( .I1(n15883), .I2(n20255), .O(n19783) );
  MUX2S U19685 ( .A(n29587), .B(n20255), .S(gray_img[1042]), .O(n19782) );
  MUX2S U19686 ( .A(n20842), .B(n20099), .S(gray_img[1018]), .O(n19428) );
  ND2S U19687 ( .I1(n15883), .I2(n20562), .O(n20564) );
  MUX2S U19688 ( .A(n20808), .B(n20562), .S(gray_img[1010]), .O(n20563) );
  AO12S U19689 ( .B1(n15883), .B2(n27829), .A1(n26221), .O(n14609) );
  AO12S U19690 ( .B1(n15935), .B2(n27081), .A1(n27073), .O(n14610) );
  AO12S U19691 ( .B1(n15883), .B2(n27065), .A1(n27057), .O(n14611) );
  AO12S U19692 ( .B1(n15883), .B2(n27261), .A1(n27187), .O(n14612) );
  MUX2S U19693 ( .A(n29587), .B(n20580), .S(gray_img[962]), .O(n19597) );
  ND2S U19694 ( .I1(n15937), .I2(n20452), .O(n18701) );
  MUX2S U19695 ( .A(n30005), .B(n20452), .S(gray_img[890]), .O(n18700) );
  ND2S U19696 ( .I1(n15937), .I2(n20559), .O(n20561) );
  MUX2S U19697 ( .A(n30005), .B(n20559), .S(gray_img[882]), .O(n20560) );
  AO12S U19698 ( .B1(n15882), .B2(n26224), .A1(n26216), .O(n14617) );
  AO12S U19699 ( .B1(n15882), .B2(n27190), .A1(n27183), .O(n14620) );
  ND2S U19700 ( .I1(n19917), .I2(n19916), .O(n14621) );
  MUX2S U19701 ( .A(n20634), .B(n20842), .S(n22988), .O(n19916) );
  MUX2S U19702 ( .A(n30005), .B(n20568), .S(gray_img[762]), .O(n19430) );
  MUX2S U19703 ( .A(n15904), .B(n20054), .S(gray_img[754]), .O(n19432) );
  ND2S U19704 ( .I1(n15937), .I2(n20365), .O(n18919) );
  MUX2S U19705 ( .A(n30005), .B(n20365), .S(gray_img[746]), .O(n18920) );
  AO12S U19706 ( .B1(n15882), .B2(n26155), .A1(n26148), .O(n14625) );
  AO12S U19707 ( .B1(n15938), .B2(n26996), .A1(n26988), .O(n14626) );
  MUX2S U19708 ( .A(n27447), .B(n26994), .S(gray_img[730]), .O(n26988) );
  AO12S U19709 ( .B1(n15882), .B2(n27009), .A1(n27001), .O(n14627) );
  AO12S U19710 ( .B1(n15882), .B2(n27243), .A1(n27130), .O(n14628) );
  ND2S U19711 ( .I1(n19882), .I2(n19881), .O(n14629) );
  ND2S U19712 ( .I1(n15937), .I2(n20623), .O(n19882) );
  MUX2S U19713 ( .A(n25928), .B(n20565), .S(gray_img[634]), .O(n19434) );
  ND2S U19714 ( .I1(n15937), .I2(n20534), .O(n20536) );
  MUX2S U19715 ( .A(n30050), .B(n20534), .S(gray_img[626]), .O(n20535) );
  ND2S U19716 ( .I1(n19852), .I2(n19851), .O(n14632) );
  ND2S U19717 ( .I1(n15937), .I2(n20274), .O(n19852) );
  MUX2S U19718 ( .A(n20274), .B(n29587), .S(n26189), .O(n19851) );
  AO12S U19719 ( .B1(n15883), .B2(n26160), .A1(n26152), .O(n14633) );
  AO12S U19720 ( .B1(n15883), .B2(n27105), .A1(n26993), .O(n14634) );
  MUX2S U19721 ( .A(n27447), .B(n27103), .S(gray_img[602]), .O(n26993) );
  AO12S U19722 ( .B1(n15882), .B2(n27013), .A1(n27006), .O(n14635) );
  MUX2S U19723 ( .A(n27447), .B(n27011), .S(gray_img[594]), .O(n27006) );
  AO12S U19724 ( .B1(n15883), .B2(n27133), .A1(n27125), .O(n14636) );
  MUX2S U19725 ( .A(n29587), .B(n20591), .S(gray_img[578]), .O(n19573) );
  ND2S U19726 ( .I1(n15937), .I2(n20472), .O(n18695) );
  MUX2S U19727 ( .A(n30056), .B(n20472), .S(gray_img[506]), .O(n18694) );
  ND2S U19728 ( .I1(n15937), .I2(n20477), .O(n18489) );
  MUX2S U19729 ( .A(n30056), .B(n20477), .S(gray_img[498]), .O(n18488) );
  ND2S U19730 ( .I1(n15937), .I2(n20480), .O(n19823) );
  MUX2S U19731 ( .A(n29597), .B(n20480), .S(gray_img[490]), .O(n19822) );
  AO12S U19732 ( .B1(n15883), .B2(n27774), .A1(n27445), .O(n14641) );
  MUX2S U19733 ( .A(n27447), .B(n27772), .S(gray_img[482]), .O(n27445) );
  AO12S U19734 ( .B1(n15883), .B2(n27352), .A1(n26756), .O(n14642) );
  AO12S U19735 ( .B1(n15883), .B2(n26747), .A1(n26744), .O(n14643) );
  MUX2S U19736 ( .A(n27447), .B(n26745), .S(gray_img[466]), .O(n26744) );
  AO12S U19737 ( .B1(n15883), .B2(n26942), .A1(n26858), .O(n14644) );
  ND2S U19738 ( .I1(n15937), .I2(n20486), .O(n18699) );
  MUX2S U19739 ( .A(n25928), .B(n20486), .S(gray_img[378]), .O(n18698) );
  ND2S U19740 ( .I1(n15883), .I2(n20522), .O(n18486) );
  MUX2S U19741 ( .A(n30050), .B(n20522), .S(gray_img[370]), .O(n18485) );
  ND2S U19742 ( .I1(n15883), .I2(n20491), .O(n19819) );
  MUX2S U19743 ( .A(n29587), .B(n20491), .S(gray_img[362]), .O(n19818) );
  AO12S U19744 ( .B1(n15883), .B2(n27449), .A1(n27440), .O(n14649) );
  MUX2S U19745 ( .A(n27447), .B(n27446), .S(gray_img[354]), .O(n27440) );
  AO12S U19746 ( .B1(n15882), .B2(n26759), .A1(n26751), .O(n14650) );
  AO12S U19747 ( .B1(n15883), .B2(n26743), .A1(n26735), .O(n14651) );
  MUX2S U19748 ( .A(n27447), .B(n26741), .S(gray_img[338]), .O(n26735) );
  AO12S U19749 ( .B1(n15935), .B2(n26861), .A1(n26853), .O(n14652) );
  ND2S U19750 ( .I1(n15883), .I2(n20496), .O(n18712) );
  MUX2S U19751 ( .A(n29597), .B(n20496), .S(gray_img[250]), .O(n18711) );
  ND2S U19752 ( .I1(n19753), .I2(n19752), .O(n14655) );
  ND2S U19753 ( .I1(n15883), .I2(n20260), .O(n19753) );
  MUX2S U19754 ( .A(n30056), .B(n20260), .S(gray_img[242]), .O(n19752) );
  ND2S U19755 ( .I1(n15883), .I2(n20620), .O(n19843) );
  MUX2S U19756 ( .A(n20842), .B(n20620), .S(gray_img[234]), .O(n19842) );
  AO12S U19757 ( .B1(n15882), .B2(n27390), .A1(n27382), .O(n14657) );
  MUX2S U19758 ( .A(n27447), .B(n27388), .S(gray_img[226]), .O(n27382) );
  AO12S U19759 ( .B1(n15882), .B2(n26726), .A1(n26706), .O(n14658) );
  AO12S U19760 ( .B1(n15882), .B2(n26841), .A1(n26719), .O(n14659) );
  AO12S U19761 ( .B1(n15882), .B2(n26883), .A1(n26876), .O(n14660) );
  ND2S U19762 ( .I1(n19903), .I2(n19902), .O(n14661) );
  ND2S U19763 ( .I1(n15883), .I2(n20631), .O(n19903) );
  MUX2S U19764 ( .A(n29587), .B(n20631), .S(gray_img[194]), .O(n19902) );
  ND2S U19765 ( .I1(n15883), .I2(n20082), .O(n18842) );
  MUX2S U19766 ( .A(n20808), .B(n20082), .S(gray_img[122]), .O(n18841) );
  ND2S U19767 ( .I1(n19757), .I2(n19756), .O(n14663) );
  ND2S U19768 ( .I1(n15883), .I2(n20499), .O(n19757) );
  MUX2S U19769 ( .A(n30056), .B(n20499), .S(gray_img[114]), .O(n19756) );
  ND2S U19770 ( .I1(n15883), .I2(n20617), .O(n19862) );
  MUX2S U19771 ( .A(n29597), .B(n20617), .S(gray_img[106]), .O(n19861) );
  AO12S U19772 ( .B1(n15882), .B2(n27545), .A1(n27387), .O(n14665) );
  MUX2S U19773 ( .A(n27447), .B(n27543), .S(gray_img[98]), .O(n27387) );
  AO12S U19774 ( .B1(n15882), .B2(n26709), .A1(n26701), .O(n14666) );
  AO12S U19775 ( .B1(n15882), .B2(n26722), .A1(n26714), .O(n14667) );
  AO12S U19776 ( .B1(n15882), .B2(n26879), .A1(n26871), .O(n14668) );
  ND2S U19777 ( .I1(n20627), .I2(n20626), .O(n14669) );
  ND2S U19778 ( .I1(n15937), .I2(n20628), .O(n20627) );
  ND2S U19779 ( .I1(n22435), .I2(n22434), .O(n15813) );
  ND3S U19780 ( .I1(n22379), .I2(n22378), .I3(n22377), .O(n22433) );
  ND2S U19781 ( .I1(n30120), .I2(n23463), .O(n23466) );
  AO12S U19782 ( .B1(n28847), .B2(n28795), .A1(n28794), .O(n14675) );
  ND2S U19783 ( .I1(n15927), .I2(n28840), .O(n28791) );
  MUX2S U19784 ( .A(n29587), .B(n28840), .S(gray_img[139]), .O(n28792) );
  ND2S U19785 ( .I1(n28727), .I2(n28226), .O(n28229) );
  OA12S U19786 ( .B1(n29843), .B2(n28730), .A1(n28227), .O(n28228) );
  MUX2S U19787 ( .A(n15904), .B(n28728), .S(gray_img[411]), .O(n28227) );
  AO12S U19788 ( .B1(n28724), .B2(n26067), .A1(n26066), .O(n13635) );
  ND2S U19789 ( .I1(n15887), .I2(n28718), .O(n26063) );
  MUX2S U19790 ( .A(n15904), .B(n28718), .S(gray_img[955]), .O(n26064) );
  AO12S U19791 ( .B1(n26096), .B2(n25922), .A1(n25921), .O(n13636) );
  ND2S U19792 ( .I1(n15927), .I2(n26090), .O(n25918) );
  MUX2S U19793 ( .A(n15904), .B(n26090), .S(gray_img[947]), .O(n25919) );
  ND2S U19794 ( .I1(n28806), .I2(n28695), .O(n28698) );
  MUX2S U19795 ( .A(n29597), .B(n28807), .S(gray_img[403]), .O(n28696) );
  AO12S U19796 ( .B1(n25619), .B2(n25597), .A1(n25596), .O(n13637) );
  ND2S U19797 ( .I1(n15887), .I2(n25612), .O(n25593) );
  MUX2S U19798 ( .A(n29566), .B(n25612), .S(gray_img[939]), .O(n25594) );
  AO12S U19799 ( .B1(n25758), .B2(n25734), .A1(n25733), .O(n13638) );
  ND2S U19800 ( .I1(n15927), .I2(n25751), .O(n25730) );
  MUX2S U19801 ( .A(n29587), .B(n25751), .S(gray_img[931]), .O(n25731) );
  AO12S U19802 ( .B1(n30128), .B2(n30055), .A1(n30054), .O(n14676) );
  ND2S U19803 ( .I1(n15925), .I2(n30121), .O(n30051) );
  MUX2S U19804 ( .A(n30050), .B(n30121), .S(gray_img[131]), .O(n30052) );
  AO12S U19805 ( .B1(n30038), .B2(n29368), .A1(n29367), .O(n14674) );
  ND2S U19806 ( .I1(n15925), .I2(n30032), .O(n29364) );
  MUX2S U19807 ( .A(n29566), .B(n30032), .S(gray_img[395]), .O(n29365) );
  MUX2S U19808 ( .A(n30056), .B(n23195), .S(gray_img[923]), .O(n23169) );
  ND2S U19809 ( .I1(n30020), .I2(n29172), .O(n29175) );
  OA12S U19810 ( .B1(n29843), .B2(n30023), .A1(n29173), .O(n29174) );
  MUX2S U19811 ( .A(n29566), .B(n30021), .S(gray_img[915]), .O(n29173) );
  AO12S U19812 ( .B1(n30109), .B2(n29985), .A1(n29984), .O(n14870) );
  ND2S U19813 ( .I1(n15925), .I2(n30103), .O(n29981) );
  MUX2S U19814 ( .A(n30056), .B(n30103), .S(gray_img[387]), .O(n29982) );
  AO12S U19815 ( .B1(n29604), .B2(n29571), .A1(n29570), .O(n13641) );
  ND2S U19816 ( .I1(n15925), .I2(n29598), .O(n29567) );
  MUX2S U19817 ( .A(n29566), .B(n29598), .S(gray_img[907]), .O(n29568) );
  AO12S U19818 ( .B1(n30098), .B2(n29471), .A1(n29470), .O(n13642) );
  ND2S U19819 ( .I1(n15927), .I2(n30092), .O(n29467) );
  MUX2S U19820 ( .A(n29587), .B(n30092), .S(gray_img[899]), .O(n29468) );
  AO12S U19821 ( .B1(n26080), .B2(n26039), .A1(n26038), .O(n13643) );
  ND2S U19822 ( .I1(n15927), .I2(n26073), .O(n26035) );
  MUX2S U19823 ( .A(n15904), .B(n26073), .S(gray_img[827]), .O(n26036) );
  AO12S U19824 ( .B1(n25936), .B2(n25891), .A1(n25890), .O(n13644) );
  MUX2S U19825 ( .A(n25928), .B(n25929), .S(gray_img[819]), .O(n25888) );
  OA12S U19826 ( .B1(n29843), .B2(n25607), .A1(n25565), .O(n25566) );
  MUX2S U19827 ( .A(n25928), .B(n25605), .S(gray_img[811]), .O(n25565) );
  AO12S U19828 ( .B1(n25750), .B2(n25709), .A1(n25708), .O(n13646) );
  ND2S U19829 ( .I1(n15927), .I2(n25744), .O(n25705) );
  MUX2S U19830 ( .A(n25928), .B(n25744), .S(gray_img[803]), .O(n25706) );
  AO12S U19831 ( .B1(n29273), .B2(n29252), .A1(n29251), .O(n13647) );
  ND2S U19832 ( .I1(n15887), .I2(n29266), .O(n29248) );
  MUX2S U19833 ( .A(n30044), .B(n29266), .S(gray_img[795]), .O(n29249) );
  AO12S U19834 ( .B1(n29192), .B2(n29151), .A1(n29150), .O(n13648) );
  ND2S U19835 ( .I1(n15925), .I2(n29186), .O(n29147) );
  MUX2S U19836 ( .A(n15904), .B(n29186), .S(gray_img[787]), .O(n29148) );
  AO12S U19837 ( .B1(n29487), .B2(n29446), .A1(n29445), .O(n13650) );
  MUX2S U19838 ( .A(n29597), .B(n29481), .S(gray_img[771]), .O(n29443) );
  ND2S U19839 ( .I1(n28247), .I2(n28191), .O(n28194) );
  OA12S U19840 ( .B1(n29843), .B2(n28250), .A1(n28192), .O(n28193) );
  MUX2S U19841 ( .A(n30005), .B(n28248), .S(gray_img[283]), .O(n28192) );
  OA12S U19842 ( .B1(n29843), .B2(n28709), .A1(n28660), .O(n28661) );
  MUX2S U19843 ( .A(n15904), .B(n28707), .S(gray_img[275]), .O(n28660) );
  AO12S U19844 ( .B1(n29381), .B2(n29334), .A1(n29333), .O(n13704) );
  ND2S U19845 ( .I1(n15927), .I2(n29374), .O(n29330) );
  MUX2S U19846 ( .A(n29587), .B(n29374), .S(gray_img[267]), .O(n29331) );
  AO12S U19847 ( .B1(n30012), .B2(n29960), .A1(n29959), .O(n13733) );
  ND2S U19848 ( .I1(n15927), .I2(n30006), .O(n29956) );
  MUX2S U19849 ( .A(n30005), .B(n30006), .S(gray_img[259]), .O(n29957) );
  AO12S U19850 ( .B1(n30087), .B2(n28834), .A1(n28833), .O(n13751) );
  ND2S U19851 ( .I1(n15927), .I2(n30081), .O(n28830) );
  MUX2S U19852 ( .A(n29566), .B(n30081), .S(gray_img[11]), .O(n28831) );
  AO12S U19853 ( .B1(n27851), .B2(n27808), .A1(n27807), .O(n13759) );
  MUX2S U19854 ( .A(n15904), .B(n27845), .S(gray_img[155]), .O(n27805) );
  AO12S U19855 ( .B1(n30076), .B2(n27319), .A1(n27318), .O(n13769) );
  ND2S U19856 ( .I1(n15927), .I2(n30070), .O(n27315) );
  MUX2S U19857 ( .A(n29566), .B(n30070), .S(gray_img[147]), .O(n27316) );
  AO12S U19858 ( .B1(n27821), .B2(n27766), .A1(n27765), .O(n13789) );
  ND2S U19859 ( .I1(n15927), .I2(n27814), .O(n27762) );
  MUX2S U19860 ( .A(n30005), .B(n27814), .S(gray_img[27]), .O(n27763) );
  AO12S U19861 ( .B1(n27378), .B2(n27344), .A1(n27343), .O(n13799) );
  ND2S U19862 ( .I1(n15927), .I2(n27371), .O(n27340) );
  MUX2S U19863 ( .A(n30005), .B(n27371), .S(gray_img[19]), .O(n27341) );
  AO12S U19864 ( .B1(n28214), .B2(n28115), .A1(n28114), .O(n13934) );
  ND2S U19865 ( .I1(n15887), .I2(n28208), .O(n28111) );
  MUX2S U19866 ( .A(n30005), .B(n28208), .S(gray_img[691]), .O(n28112) );
  AO12S U19867 ( .B1(n28607), .B2(n28446), .A1(n28445), .O(n13941) );
  ND2S U19868 ( .I1(n15927), .I2(n28601), .O(n28442) );
  MUX2S U19869 ( .A(n15904), .B(n28601), .S(gray_img[683]), .O(n28443) );
  AO12S U19870 ( .B1(n28588), .B2(n28552), .A1(n28551), .O(n13948) );
  ND2S U19871 ( .I1(n15927), .I2(n28581), .O(n28548) );
  MUX2S U19872 ( .A(n30056), .B(n28581), .S(gray_img[675]), .O(n28549) );
  AO12S U19873 ( .B1(n29350), .B2(n28909), .A1(n28908), .O(n13956) );
  ND2S U19874 ( .I1(n15925), .I2(n29344), .O(n28905) );
  MUX2S U19875 ( .A(n29597), .B(n29344), .S(gray_img[667]), .O(n28906) );
  AO12S U19876 ( .B1(n29040), .B2(n29003), .A1(n29002), .O(n13964) );
  ND2S U19877 ( .I1(n15887), .I2(n29033), .O(n28999) );
  MUX2S U19878 ( .A(n29566), .B(n29033), .S(gray_img[659]), .O(n29000) );
  AO12S U19879 ( .B1(n29904), .B2(n29873), .A1(n29872), .O(n13973) );
  ND2S U19880 ( .I1(n15927), .I2(n29898), .O(n29869) );
  MUX2S U19881 ( .A(n30044), .B(n29898), .S(gray_img[651]), .O(n29870) );
  ND2S U19882 ( .I1(n29993), .I2(n29696), .O(n29699) );
  OA12S U19883 ( .B1(n29843), .B2(n29996), .A1(n29697), .O(n29698) );
  MUX2S U19884 ( .A(n15904), .B(n29994), .S(gray_img[643]), .O(n29697) );
  ND2S U19885 ( .I1(n23492), .I2(n23345), .O(n23348) );
  MUX2S U19886 ( .A(n30044), .B(n23493), .S(gray_img[571]), .O(n23346) );
  AO12S U19887 ( .B1(n28128), .B2(n28084), .A1(n28083), .O(n14016) );
  ND2S U19888 ( .I1(n15927), .I2(n28121), .O(n28080) );
  MUX2S U19889 ( .A(n30005), .B(n28121), .S(gray_img[563]), .O(n28081) );
  AO12S U19890 ( .B1(n28459), .B2(n28415), .A1(n28414), .O(n14025) );
  ND2S U19891 ( .I1(n15927), .I2(n28452), .O(n28411) );
  MUX2S U19892 ( .A(n29032), .B(n28452), .S(gray_img[555]), .O(n28412) );
  ND2S U19893 ( .I1(n28671), .I2(n28571), .O(n28574) );
  OA12S U19894 ( .B1(n29843), .B2(n28674), .A1(n28572), .O(n28573) );
  MUX2S U19895 ( .A(n15904), .B(n28672), .S(gray_img[547]), .O(n28572) );
  AO12S U19896 ( .B1(n28950), .B2(n28929), .A1(n28928), .O(n14043) );
  ND2S U19897 ( .I1(n15927), .I2(n28943), .O(n28925) );
  MUX2S U19898 ( .A(n30056), .B(n28943), .S(gray_img[539]), .O(n28926) );
  ND2S U19899 ( .I1(n29043), .I2(n29027), .O(n29030) );
  MUX2S U19900 ( .A(n30056), .B(n29044), .S(gray_img[531]), .O(n29028) );
  OA12S U19901 ( .B1(n29843), .B2(n29883), .A1(n29842), .O(n29844) );
  MUX2S U19902 ( .A(n30005), .B(n29881), .S(gray_img[523]), .O(n29842) );
  OA12S U19903 ( .B1(n29843), .B2(n29742), .A1(n29722), .O(n29723) );
  MUX2S U19904 ( .A(n15904), .B(n29740), .S(gray_img[515]), .O(n29722) );
  AO12S U19905 ( .B1(n26473), .B2(n26431), .A1(n26430), .O(n14095) );
  ND2S U19906 ( .I1(n15927), .I2(n26466), .O(n26427) );
  MUX2S U19907 ( .A(n15904), .B(n26466), .S(gray_img[443]), .O(n26428) );
  AO12S U19908 ( .B1(n27840), .B2(n26286), .A1(n26285), .O(n14104) );
  ND2S U19909 ( .I1(n15887), .I2(n27834), .O(n26282) );
  MUX2S U19910 ( .A(n30056), .B(n27834), .S(gray_img[435]), .O(n26283) );
  ND2S U19911 ( .I1(n23121), .I2(n23100), .O(n23103) );
  MUX2S U19912 ( .A(n29597), .B(n25151), .S(gray_img[427]), .O(n23101) );
  OA12S U19913 ( .B1(n29843), .B2(n27224), .A1(n27212), .O(n27215) );
  ND2S U19914 ( .I1(n27226), .I2(n27213), .O(n27214) );
  MUX2S U19915 ( .A(n30050), .B(n27222), .S(gray_img[419]), .O(n27212) );
  AO12S U19916 ( .B1(n26489), .B2(n26460), .A1(n26459), .O(n14139) );
  ND2S U19917 ( .I1(n15927), .I2(n26483), .O(n26456) );
  MUX2S U19918 ( .A(n30044), .B(n26483), .S(gray_img[315]), .O(n26457) );
  ND2S U19919 ( .I1(n26327), .I2(n26308), .O(n26309) );
  OA12S U19920 ( .B1(n29843), .B2(n26324), .A1(n26307), .O(n26310) );
  MUX2S U19921 ( .A(n15904), .B(n26322), .S(gray_img[307]), .O(n26307) );
  AO12S U19922 ( .B1(n27121), .B2(n27097), .A1(n27096), .O(n14157) );
  ND2S U19923 ( .I1(n15927), .I2(n27114), .O(n27093) );
  MUX2S U19924 ( .A(n29597), .B(n27114), .S(gray_img[299]), .O(n27094) );
  OA12S U19925 ( .B1(n29843), .B2(n27254), .A1(n27232), .O(n27233) );
  ND2S U19926 ( .I1(n27251), .I2(n27231), .O(n27234) );
  MUX2S U19927 ( .A(n29566), .B(n27252), .S(gray_img[291]), .O(n27232) );
  AO12S U19928 ( .B1(n27692), .B2(n27651), .A1(n27650), .O(n14183) );
  ND2S U19929 ( .I1(n15925), .I2(n27685), .O(n27647) );
  MUX2S U19930 ( .A(n30044), .B(n27685), .S(gray_img[187]), .O(n27648) );
  AO12S U19931 ( .B1(n27785), .B2(n27506), .A1(n27505), .O(n14192) );
  ND2S U19932 ( .I1(n15927), .I2(n27779), .O(n27502) );
  MUX2S U19933 ( .A(n29587), .B(n27779), .S(gray_img[179]), .O(n27503) );
  OA12S U19934 ( .B1(n29843), .B2(n27358), .A1(n26814), .O(n26815) );
  MUX2S U19935 ( .A(n30044), .B(n27356), .S(gray_img[171]), .O(n26814) );
  AO12S U19936 ( .B1(n26939), .B2(n26918), .A1(n26917), .O(n14210) );
  ND2S U19937 ( .I1(n15887), .I2(n26932), .O(n26914) );
  MUX2S U19938 ( .A(n29032), .B(n26932), .S(gray_img[163]), .O(n26915) );
  AO12S U19939 ( .B1(n27708), .B2(n27679), .A1(n27678), .O(n14227) );
  MUX2S U19940 ( .A(n30056), .B(n27702), .S(gray_img[59]), .O(n27676) );
  AO12S U19941 ( .B1(n27556), .B2(n27532), .A1(n27531), .O(n14236) );
  ND2S U19942 ( .I1(n15927), .I2(n27550), .O(n27528) );
  MUX2S U19943 ( .A(n29032), .B(n27550), .S(gray_img[51]), .O(n27529) );
  ND2S U19944 ( .I1(n15887), .I2(n26842), .O(n16066) );
  AO12S U19945 ( .B1(n26931), .B2(n26898), .A1(n26897), .O(n14254) );
  ND2S U19946 ( .I1(n15927), .I2(n26924), .O(n26894) );
  MUX2S U19947 ( .A(n30044), .B(n26924), .S(gray_img[35]), .O(n26895) );
  ND2S U19948 ( .I1(n28136), .I2(n27944), .O(n27947) );
  OA12S U19949 ( .B1(n29843), .B2(n28139), .A1(n27945), .O(n27946) );
  MUX2S U19950 ( .A(n30005), .B(n28137), .S(gray_img[699]), .O(n27945) );
  ND2S U19951 ( .I1(n15880), .I2(n25942), .O(n18583) );
  AO12S U19952 ( .B1(n15927), .B2(n25836), .A1(n25828), .O(n14681) );
  MUX2S U19953 ( .A(n15889), .B(n25834), .S(gray_img[2019]), .O(n25828) );
  AO12S U19954 ( .B1(n15925), .B2(n25473), .A1(n25464), .O(n14682) );
  MUX2S U19955 ( .A(n28534), .B(n25471), .S(gray_img[2011]), .O(n25464) );
  AO12S U19956 ( .B1(n15927), .B2(n25761), .A1(n25456), .O(n14683) );
  MUX2S U19957 ( .A(n28534), .B(n25759), .S(gray_img[2003]), .O(n25456) );
  AO12S U19958 ( .B1(n15927), .B2(n28803), .A1(n25627), .O(n14684) );
  MUX2S U19959 ( .A(n15889), .B(n28801), .S(gray_img[1995]), .O(n25627) );
  ND2S U19960 ( .I1(n15880), .I2(n20209), .O(n18949) );
  ND2S U19961 ( .I1(n15881), .I2(n20746), .O(n20748) );
  MUX2S U19962 ( .A(n29566), .B(n20746), .S(gray_img[1979]), .O(n20747) );
  ND2S U19963 ( .I1(n15881), .I2(n20849), .O(n20850) );
  MUX2S U19964 ( .A(n29597), .B(n20849), .S(gray_img[1971]), .O(n20851) );
  MUX2S U19965 ( .A(n29566), .B(n19970), .S(gray_img[1947]), .O(n19541) );
  MUX2S U19966 ( .A(n30050), .B(n20389), .S(gray_img[1939]), .O(n19575) );
  MUX2S U19967 ( .A(n20830), .B(n20424), .S(gray_img[1931]), .O(n19524) );
  MUX2S U19968 ( .A(n20842), .B(n20373), .S(gray_img[1923]), .O(n19559) );
  ND2S U19969 ( .I1(n15881), .I2(n20430), .O(n18788) );
  MUX2S U19970 ( .A(n30044), .B(n20430), .S(gray_img[1915]), .O(n18787) );
  ND2S U19971 ( .I1(n15881), .I2(n20063), .O(n18497) );
  MUX2S U19972 ( .A(n29566), .B(n20063), .S(gray_img[1907]), .O(n18496) );
  MUX2S U19973 ( .A(n30056), .B(n20544), .S(gray_img[1899]), .O(n19438) );
  AO12S U19974 ( .B1(n15926), .B2(n25832), .A1(n25823), .O(n14697) );
  MUX2S U19975 ( .A(n27447), .B(n25830), .S(gray_img[1891]), .O(n25823) );
  AO12S U19976 ( .B1(n15927), .B2(n25477), .A1(n25469), .O(n14698) );
  AO12S U19977 ( .B1(n15925), .B2(n25460), .A1(n25452), .O(n14699) );
  AO12S U19978 ( .B1(n15887), .B2(n25631), .A1(n25622), .O(n14700) );
  MUX2S U19979 ( .A(n15889), .B(n25629), .S(gray_img[1867]), .O(n25622) );
  MUX2S U19980 ( .A(n20842), .B(n20504), .S(gray_img[1859]), .O(n19442) );
  ND2S U19981 ( .I1(n15881), .I2(n20740), .O(n20742) );
  MUX2S U19982 ( .A(n29566), .B(n20740), .S(gray_img[1851]), .O(n20741) );
  ND2S U19983 ( .I1(n15881), .I2(n20862), .O(n20860) );
  MUX2S U19984 ( .A(n29597), .B(n20862), .S(gray_img[1843]), .O(n20861) );
  ND2S U19985 ( .I1(n15881), .I2(n20142), .O(n18766) );
  ND2S U19986 ( .I1(n15881), .I2(n20156), .O(n18472) );
  MUX2S U19987 ( .A(n29587), .B(n20296), .S(gray_img[1819]), .O(n19599) );
  MUX2S U19988 ( .A(n29597), .B(n20354), .S(gray_img[1811]), .O(n20345) );
  MUX2S U19989 ( .A(n20830), .B(n20319), .S(gray_img[1803]), .O(n19450) );
  MUX2S U19990 ( .A(n29587), .B(n20376), .S(gray_img[1795]), .O(n19587) );
  ND2S U19991 ( .I1(n15881), .I2(n20547), .O(n18794) );
  MUX2S U19992 ( .A(n29566), .B(n20547), .S(gray_img[1787]), .O(n18793) );
  ND2S U19993 ( .I1(n15881), .I2(n20541), .O(n18491) );
  MUX2S U19994 ( .A(n29587), .B(n20541), .S(gray_img[1779]), .O(n18490) );
  MUX2S U19995 ( .A(n29597), .B(n20449), .S(gray_img[1771]), .O(n19456) );
  AO12S U19996 ( .B1(n15887), .B2(n25778), .A1(n25769), .O(n14713) );
  MUX2S U19997 ( .A(n27447), .B(n25776), .S(gray_img[1763]), .O(n25769) );
  AO12S U19998 ( .B1(n15887), .B2(n25510), .A1(n25501), .O(n14714) );
  AO12S U19999 ( .B1(n15887), .B2(n25498), .A1(n25490), .O(n14715) );
  MUX2S U20000 ( .A(n28534), .B(n25496), .S(gray_img[1747]), .O(n25490) );
  AO12S U20001 ( .B1(n15880), .B2(n25649), .A1(n25640), .O(n14716) );
  MUX2S U20002 ( .A(n15889), .B(n25647), .S(gray_img[1739]), .O(n25640) );
  MUX2S U20003 ( .A(n30056), .B(n19955), .S(gray_img[1731]), .O(n19464) );
  ND2S U20004 ( .I1(n15881), .I2(n20737), .O(n20713) );
  MUX2S U20005 ( .A(n30056), .B(n20737), .S(gray_img[1723]), .O(n20712) );
  ND2S U20006 ( .I1(n15881), .I2(n20846), .O(n20847) );
  MUX2S U20007 ( .A(n30050), .B(n20846), .S(gray_img[1715]), .O(n20848) );
  ND2S U20008 ( .I1(n15881), .I2(n20827), .O(n20794) );
  MUX2S U20009 ( .A(n30050), .B(n20827), .S(gray_img[1707]), .O(n20795) );
  ND2S U20010 ( .I1(n15881), .I2(n20787), .O(n19656) );
  MUX2S U20011 ( .A(n30056), .B(n20787), .S(gray_img[1699]), .O(n19657) );
  ND2S U20012 ( .I1(n15881), .I2(n20599), .O(n20600) );
  MUX2S U20013 ( .A(n29597), .B(n20599), .S(gray_img[1691]), .O(n20601) );
  ND2S U20014 ( .I1(n15881), .I2(n20605), .O(n20606) );
  MUX2S U20015 ( .A(n29566), .B(n20605), .S(gray_img[1683]), .O(n20607) );
  ND2S U20016 ( .I1(n15881), .I2(n20531), .O(n20508) );
  MUX2S U20017 ( .A(n29597), .B(n20531), .S(gray_img[1675]), .O(n20507) );
  ND2S U20018 ( .I1(n15881), .I2(n20583), .O(n20576) );
  MUX2S U20019 ( .A(n29587), .B(n20583), .S(gray_img[1667]), .O(n20577) );
  ND2S U20020 ( .I1(n15881), .I2(n20509), .O(n18798) );
  MUX2S U20021 ( .A(n29597), .B(n20509), .S(gray_img[1659]), .O(n18797) );
  ND2S U20022 ( .I1(n15881), .I2(n20525), .O(n18494) );
  MUX2S U20023 ( .A(n29587), .B(n20525), .S(gray_img[1651]), .O(n18493) );
  MUX2S U20024 ( .A(n29597), .B(n20463), .S(gray_img[1643]), .O(n19466) );
  AO12S U20025 ( .B1(n15881), .B2(n25899), .A1(n25774), .O(n14729) );
  MUX2S U20026 ( .A(n15889), .B(n25897), .S(gray_img[1635]), .O(n25774) );
  AO12S U20027 ( .B1(n15881), .B2(n25576), .A1(n25506), .O(n14730) );
  MUX2S U20028 ( .A(n27447), .B(n25574), .S(gray_img[1627]), .O(n25506) );
  AO12S U20029 ( .B1(n15887), .B2(n25494), .A1(n25485), .O(n14731) );
  MUX2S U20030 ( .A(n28534), .B(n25492), .S(gray_img[1619]), .O(n25485) );
  AO12S U20031 ( .B1(n15880), .B2(n25653), .A1(n25645), .O(n14732) );
  MUX2S U20032 ( .A(n30050), .B(n20528), .S(gray_img[1603]), .O(n19478) );
  ND2S U20033 ( .I1(n15881), .I2(n20731), .O(n20733) );
  MUX2S U20034 ( .A(n30050), .B(n20731), .S(gray_img[1595]), .O(n20732) );
  ND2S U20035 ( .I1(n15881), .I2(n20839), .O(n20840) );
  MUX2S U20036 ( .A(n30056), .B(n20839), .S(gray_img[1587]), .O(n20841) );
  ND2S U20037 ( .I1(n15881), .I2(n20395), .O(n19662) );
  MUX2S U20038 ( .A(n30050), .B(n20395), .S(gray_img[1579]), .O(n19663) );
  ND2S U20039 ( .I1(n15880), .I2(n20824), .O(n20825) );
  MUX2S U20040 ( .A(n30056), .B(n20824), .S(gray_img[1571]), .O(n20826) );
  ND2S U20041 ( .I1(n15880), .I2(n20596), .O(n20597) );
  MUX2S U20042 ( .A(n29566), .B(n20596), .S(gray_img[1563]), .O(n20598) );
  ND2S U20043 ( .I1(n15880), .I2(n20602), .O(n20594) );
  MUX2S U20044 ( .A(n29597), .B(n20602), .S(gray_img[1555]), .O(n20595) );
  ND2S U20045 ( .I1(n15880), .I2(n20550), .O(n20552) );
  MUX2S U20046 ( .A(n29566), .B(n20550), .S(gray_img[1547]), .O(n20551) );
  ND2S U20047 ( .I1(n15880), .I2(n20881), .O(n20867) );
  MUX2S U20048 ( .A(n29597), .B(n20881), .S(gray_img[1539]), .O(n20868) );
  ND2S U20049 ( .I1(n15880), .I2(n20556), .O(n20558) );
  MUX2S U20050 ( .A(n30044), .B(n20556), .S(gray_img[1531]), .O(n20557) );
  ND2S U20051 ( .I1(n15880), .I2(n20512), .O(n20514) );
  MUX2S U20052 ( .A(n20830), .B(n20512), .S(gray_img[1523]), .O(n20513) );
  ND2S U20053 ( .I1(n15880), .I2(n20440), .O(n19637) );
  MUX2S U20054 ( .A(n30056), .B(n20440), .S(gray_img[1515]), .O(n19636) );
  AO12S U20055 ( .B1(n15880), .B2(n27971), .A1(n27963), .O(n14745) );
  MUX2S U20056 ( .A(n28534), .B(n27969), .S(gray_img[1507]), .O(n27963) );
  AO12S U20057 ( .B1(n15926), .B2(n28355), .A1(n28346), .O(n14746) );
  AO12S U20058 ( .B1(n15880), .B2(n28342), .A1(n28333), .O(n14747) );
  MUX2S U20059 ( .A(n27447), .B(n28340), .S(gray_img[1491]), .O(n28333) );
  AO12S U20060 ( .B1(n15887), .B2(n28560), .A1(n28531), .O(n14748) );
  ND2S U20061 ( .I1(n15880), .I2(n20684), .O(n20686) );
  MUX2S U20062 ( .A(n30056), .B(n20684), .S(gray_img[1475]), .O(n20685) );
  ND2S U20063 ( .I1(n15880), .I2(n20709), .O(n20675) );
  ND2S U20064 ( .I1(n15880), .I2(n20821), .O(n20817) );
  MUX2S U20065 ( .A(n30044), .B(n20821), .S(gray_img[1459]), .O(n20818) );
  ND2S U20066 ( .I1(n15880), .I2(n20814), .O(n20815) );
  MUX2S U20067 ( .A(n29566), .B(n20814), .S(gray_img[1451]), .O(n20816) );
  ND2S U20068 ( .I1(n15880), .I2(n20811), .O(n20812) );
  ND2S U20069 ( .I1(n15880), .I2(n20293), .O(n18629) );
  MUX2S U20070 ( .A(n30056), .B(n20293), .S(gray_img[1435]), .O(n18630) );
  MUX2S U20071 ( .A(n20842), .B(n20193), .S(gray_img[1427]), .O(n19589) );
  ND2S U20072 ( .I1(n15880), .I2(n20035), .O(n18726) );
  MUX2S U20073 ( .A(n20842), .B(n20035), .S(gray_img[1419]), .O(n18725) );
  ND2S U20074 ( .I1(n15880), .I2(n20359), .O(n18868) );
  ND2S U20075 ( .I1(n15880), .I2(n20571), .O(n20573) );
  MUX2S U20076 ( .A(n30056), .B(n20571), .S(gray_img[1403]), .O(n20572) );
  ND2S U20077 ( .I1(n15880), .I2(n20517), .O(n20519) );
  MUX2S U20078 ( .A(n20808), .B(n20517), .S(gray_img[1395]), .O(n20518) );
  ND2S U20079 ( .I1(n15880), .I2(n20722), .O(n20706) );
  MUX2S U20080 ( .A(n30056), .B(n20722), .S(gray_img[1387]), .O(n20705) );
  AO12S U20081 ( .B1(n15927), .B2(n28203), .A1(n27967), .O(n14761) );
  MUX2S U20082 ( .A(n28534), .B(n28201), .S(gray_img[1379]), .O(n27967) );
  AO12S U20083 ( .B1(n15926), .B2(n28359), .A1(n28351), .O(n14762) );
  AO12S U20084 ( .B1(n15880), .B2(n28596), .A1(n28338), .O(n14763) );
  AO12S U20085 ( .B1(n15881), .B2(n28536), .A1(n28525), .O(n14764) );
  MUX2S U20086 ( .A(n28534), .B(n28533), .S(gray_img[1355]), .O(n28525) );
  ND2S U20087 ( .I1(n15880), .I2(n20734), .O(n20699) );
  MUX2S U20088 ( .A(n30044), .B(n20734), .S(gray_img[1347]), .O(n20698) );
  ND2S U20089 ( .I1(n15926), .I2(n20695), .O(n20697) );
  MUX2S U20090 ( .A(n30044), .B(n20695), .S(gray_img[1339]), .O(n20696) );
  ND2S U20091 ( .I1(n15926), .I2(n20833), .O(n20806) );
  MUX2S U20092 ( .A(n30044), .B(n20833), .S(gray_img[1331]), .O(n20807) );
  ND2S U20093 ( .I1(n15926), .I2(n20836), .O(n20804) );
  MUX2S U20094 ( .A(n29566), .B(n20836), .S(gray_img[1323]), .O(n20805) );
  ND2S U20095 ( .I1(n15926), .I2(n20843), .O(n20800) );
  MUX2S U20096 ( .A(n30056), .B(n20843), .S(gray_img[1315]), .O(n20801) );
  MUX2S U20097 ( .A(n29566), .B(n20362), .S(gray_img[1299]), .O(n19583) );
  ND2S U20098 ( .I1(n15926), .I2(n20427), .O(n18732) );
  MUX2S U20099 ( .A(n20842), .B(n20427), .S(gray_img[1291]), .O(n18731) );
  ND2S U20100 ( .I1(n15926), .I2(n20392), .O(n18872) );
  MUX2S U20101 ( .A(n29587), .B(n20392), .S(gray_img[1283]), .O(n18873) );
  ND2S U20102 ( .I1(n15926), .I2(n20655), .O(n20648) );
  MUX2S U20103 ( .A(n20808), .B(n20655), .S(gray_img[1275]), .O(n20647) );
  ND2S U20104 ( .I1(n15926), .I2(n20725), .O(n20692) );
  MUX2S U20105 ( .A(n20808), .B(n20725), .S(gray_img[1267]), .O(n20691) );
  ND2S U20106 ( .I1(n15926), .I2(n20719), .O(n20652) );
  MUX2S U20107 ( .A(n30050), .B(n20719), .S(gray_img[1259]), .O(n20651) );
  AO12S U20108 ( .B1(n15881), .B2(n28031), .A1(n28026), .O(n14777) );
  AO12S U20109 ( .B1(n15881), .B2(n28288), .A1(n28280), .O(n14778) );
  AO12S U20110 ( .B1(n15887), .B2(n28271), .A1(n28262), .O(n14779) );
  AO12S U20111 ( .B1(n15881), .B2(n28475), .A1(n28468), .O(n14780) );
  ND2S U20112 ( .I1(n15926), .I2(n20702), .O(n20640) );
  MUX2S U20113 ( .A(n29587), .B(n20702), .S(gray_img[1219]), .O(n20639) );
  ND2S U20114 ( .I1(n20754), .I2(n20753), .O(n14782) );
  ND2S U20115 ( .I1(n15880), .I2(n20757), .O(n20754) );
  MUX2S U20116 ( .A(n30044), .B(n20757), .S(gray_img[1211]), .O(n20753) );
  ND2S U20117 ( .I1(n15927), .I2(n20857), .O(n20785) );
  MUX2S U20118 ( .A(n30044), .B(n20857), .S(gray_img[1203]), .O(n20786) );
  ND2S U20119 ( .I1(n15925), .I2(n20435), .O(n19679) );
  MUX2S U20120 ( .A(n29587), .B(n20435), .S(gray_img[1195]), .O(n19678) );
  ND2S U20121 ( .I1(n15880), .I2(n20379), .O(n18505) );
  MUX2S U20122 ( .A(n29566), .B(n20379), .S(gray_img[1187]), .O(n18506) );
  ND2S U20123 ( .I1(n15927), .I2(n20159), .O(n18635) );
  MUX2S U20124 ( .A(n29597), .B(n20159), .S(gray_img[1179]), .O(n18636) );
  ND2S U20125 ( .I1(n15927), .I2(n20316), .O(n19771) );
  MUX2S U20126 ( .A(n29597), .B(n20316), .S(gray_img[1171]), .O(n19770) );
  ND2S U20127 ( .I1(n15927), .I2(n20553), .O(n20555) );
  MUX2S U20128 ( .A(n29597), .B(n20553), .S(gray_img[1163]), .O(n20554) );
  MUX2S U20129 ( .A(n29597), .B(n20240), .S(gray_img[1155]), .O(n19706) );
  ND2S U20130 ( .I1(n15927), .I2(n20716), .O(n20646) );
  MUX2S U20131 ( .A(n30050), .B(n20716), .S(gray_img[1147]), .O(n20645) );
  ND2S U20132 ( .I1(n15927), .I2(n20124), .O(n19633) );
  MUX2S U20133 ( .A(n20808), .B(n20124), .S(gray_img[1139]), .O(n19632) );
  ND2S U20134 ( .I1(n15880), .I2(n20728), .O(n20667) );
  MUX2S U20135 ( .A(n30044), .B(n20728), .S(gray_img[1131]), .O(n20666) );
  AO12S U20136 ( .B1(n15887), .B2(n28092), .A1(n28021), .O(n14793) );
  MUX2S U20137 ( .A(n28534), .B(n28090), .S(gray_img[1123]), .O(n28021) );
  AO12S U20138 ( .B1(n15887), .B2(n28284), .A1(n28275), .O(n14794) );
  AO12S U20139 ( .B1(n15887), .B2(n28423), .A1(n28267), .O(n14795) );
  AO12S U20140 ( .B1(n15887), .B2(n28480), .A1(n28471), .O(n14796) );
  ND2S U20141 ( .I1(n15881), .I2(n20743), .O(n20669) );
  MUX2S U20142 ( .A(n30050), .B(n20743), .S(gray_img[1091]), .O(n20668) );
  ND2S U20143 ( .I1(n20762), .I2(n20761), .O(n14798) );
  ND2S U20144 ( .I1(n15926), .I2(n20760), .O(n20762) );
  MUX2S U20145 ( .A(n30056), .B(n20760), .S(gray_img[1083]), .O(n20761) );
  ND2S U20146 ( .I1(n15881), .I2(n20854), .O(n20781) );
  MUX2S U20147 ( .A(n30044), .B(n20854), .S(gray_img[1075]), .O(n20782) );
  ND2S U20148 ( .I1(n15926), .I2(n20611), .O(n19683) );
  MUX2S U20149 ( .A(n29566), .B(n20611), .S(gray_img[1067]), .O(n19682) );
  ND2S U20150 ( .I1(n15880), .I2(n20368), .O(n18514) );
  MUX2S U20151 ( .A(n29597), .B(n20368), .S(gray_img[1059]), .O(n18515) );
  MUX2S U20152 ( .A(n29587), .B(n20184), .S(gray_img[1051]), .O(n19547) );
  ND2S U20153 ( .I1(n19787), .I2(n19786), .O(n14803) );
  ND2S U20154 ( .I1(n15881), .I2(n20255), .O(n19787) );
  MUX2S U20155 ( .A(n29566), .B(n20255), .S(gray_img[1043]), .O(n19786) );
  MUX2S U20156 ( .A(n29587), .B(n20235), .S(gray_img[1035]), .O(n19644) );
  MUX2S U20157 ( .A(n15904), .B(n20099), .S(gray_img[1019]), .O(n19488) );
  ND2S U20158 ( .I1(n15880), .I2(n20562), .O(n20540) );
  MUX2S U20159 ( .A(n20830), .B(n20562), .S(gray_img[1011]), .O(n20539) );
  AO12S U20160 ( .B1(n15925), .B2(n27829), .A1(n26220), .O(n14809) );
  MUX2S U20161 ( .A(n15889), .B(n27827), .S(gray_img[995]), .O(n26220) );
  AO12S U20162 ( .B1(n15887), .B2(n27081), .A1(n27072), .O(n14810) );
  AO12S U20163 ( .B1(n15887), .B2(n27065), .A1(n27056), .O(n14811) );
  AO12S U20164 ( .B1(n15887), .B2(n27261), .A1(n27186), .O(n14812) );
  ND2S U20165 ( .I1(n15880), .I2(n20580), .O(n18943) );
  MUX2S U20166 ( .A(n29587), .B(n20580), .S(gray_img[963]), .O(n18944) );
  ND2S U20167 ( .I1(n15881), .I2(n20452), .O(n18697) );
  MUX2S U20168 ( .A(n30005), .B(n20452), .S(gray_img[891]), .O(n18696) );
  ND2S U20169 ( .I1(n15880), .I2(n20559), .O(n20538) );
  MUX2S U20170 ( .A(n30005), .B(n20559), .S(gray_img[883]), .O(n20537) );
  AO12S U20171 ( .B1(n15927), .B2(n26224), .A1(n26215), .O(n14817) );
  MUX2S U20172 ( .A(n27447), .B(n26222), .S(gray_img[867]), .O(n26215) );
  AO12S U20173 ( .B1(n15880), .B2(n30065), .A1(n27077), .O(n14818) );
  AO12S U20174 ( .B1(n15880), .B2(n27069), .A1(n27061), .O(n14819) );
  AO12S U20175 ( .B1(n15880), .B2(n27190), .A1(n27182), .O(n14820) );
  ND2S U20176 ( .I1(n19919), .I2(n19918), .O(n14821) );
  MUX2S U20177 ( .A(n20634), .B(n20808), .S(n22986), .O(n19918) );
  MUX2S U20178 ( .A(n25928), .B(n20568), .S(gray_img[763]), .O(n19494) );
  MUX2S U20179 ( .A(n30005), .B(n20054), .S(gray_img[755]), .O(n19496) );
  AO12S U20180 ( .B1(n15925), .B2(n26155), .A1(n26147), .O(n14825) );
  AO12S U20181 ( .B1(n15925), .B2(n26996), .A1(n26987), .O(n14826) );
  AO12S U20182 ( .B1(n15880), .B2(n27009), .A1(n27000), .O(n14827) );
  AO12S U20183 ( .B1(n15880), .B2(n27243), .A1(n27129), .O(n14828) );
  ND2S U20184 ( .I1(n19869), .I2(n19868), .O(n14829) );
  MUX2S U20185 ( .A(n29597), .B(n20623), .S(gray_img[707]), .O(n19868) );
  MUX2S U20186 ( .A(n30005), .B(n20565), .S(gray_img[635]), .O(n19498) );
  ND2S U20187 ( .I1(n15925), .I2(n20534), .O(n20516) );
  MUX2S U20188 ( .A(n30050), .B(n20534), .S(gray_img[627]), .O(n20515) );
  ND2S U20189 ( .I1(n19850), .I2(n19849), .O(n14832) );
  ND2S U20190 ( .I1(n15880), .I2(n20274), .O(n19850) );
  MUX2S U20191 ( .A(n20274), .B(n20830), .S(n26187), .O(n19849) );
  AO12S U20192 ( .B1(n15925), .B2(n26160), .A1(n26151), .O(n14833) );
  AO12S U20193 ( .B1(n15927), .B2(n27105), .A1(n26992), .O(n14834) );
  MUX2S U20194 ( .A(n15889), .B(n27103), .S(gray_img[603]), .O(n26992) );
  AO12S U20195 ( .B1(n15927), .B2(n27013), .A1(n27005), .O(n14835) );
  MUX2S U20196 ( .A(n27447), .B(n27011), .S(gray_img[595]), .O(n27005) );
  AO12S U20197 ( .B1(n15927), .B2(n27133), .A1(n27124), .O(n14836) );
  ND2S U20198 ( .I1(n15925), .I2(n20591), .O(n18941) );
  MUX2S U20199 ( .A(n29587), .B(n20591), .S(gray_img[579]), .O(n18942) );
  MUX2S U20200 ( .A(n30044), .B(n20477), .S(gray_img[499]), .O(n19508) );
  ND2S U20201 ( .I1(n15927), .I2(n20480), .O(n19821) );
  MUX2S U20202 ( .A(n29566), .B(n20480), .S(gray_img[491]), .O(n19820) );
  AO12S U20203 ( .B1(n15927), .B2(n27774), .A1(n27444), .O(n14841) );
  MUX2S U20204 ( .A(n27447), .B(n27772), .S(gray_img[483]), .O(n27444) );
  AO12S U20205 ( .B1(n15927), .B2(n27352), .A1(n26755), .O(n14842) );
  AO12S U20206 ( .B1(n15927), .B2(n26747), .A1(n26738), .O(n14843) );
  MUX2S U20207 ( .A(n27447), .B(n26745), .S(gray_img[467]), .O(n26738) );
  AO12S U20208 ( .B1(n15927), .B2(n26942), .A1(n26857), .O(n14844) );
  ND2S U20209 ( .I1(n19888), .I2(n19887), .O(n14845) );
  ND2S U20210 ( .I1(n15880), .I2(n20483), .O(n19888) );
  MUX2S U20211 ( .A(n30044), .B(n20486), .S(gray_img[379]), .O(n19510) );
  ND2S U20212 ( .I1(n15880), .I2(n20522), .O(n20524) );
  MUX2S U20213 ( .A(n20842), .B(n20522), .S(gray_img[371]), .O(n20523) );
  ND2S U20214 ( .I1(n15880), .I2(n20491), .O(n19817) );
  MUX2S U20215 ( .A(n29566), .B(n20491), .S(gray_img[363]), .O(n19816) );
  AO12S U20216 ( .B1(n15925), .B2(n27449), .A1(n27439), .O(n14849) );
  MUX2S U20217 ( .A(n27447), .B(n27446), .S(gray_img[355]), .O(n27439) );
  AO12S U20218 ( .B1(n15927), .B2(n26759), .A1(n26750), .O(n14850) );
  AO12S U20219 ( .B1(n15927), .B2(n26743), .A1(n26734), .O(n14851) );
  MUX2S U20220 ( .A(n28534), .B(n26741), .S(gray_img[339]), .O(n26734) );
  AO12S U20221 ( .B1(n15927), .B2(n26861), .A1(n26852), .O(n14852) );
  MUX2S U20222 ( .A(n29587), .B(n20496), .S(gray_img[251]), .O(n19512) );
  ND2S U20223 ( .I1(n19749), .I2(n19748), .O(n14855) );
  ND2S U20224 ( .I1(n15927), .I2(n20260), .O(n19749) );
  MUX2S U20225 ( .A(n30044), .B(n20260), .S(gray_img[243]), .O(n19748) );
  MUX2S U20226 ( .A(n29587), .B(n20620), .S(gray_img[235]), .O(n19831) );
  AO12S U20227 ( .B1(n15925), .B2(n27390), .A1(n27381), .O(n14857) );
  MUX2S U20228 ( .A(n27447), .B(n27388), .S(gray_img[227]), .O(n27381) );
  AO12S U20229 ( .B1(n15927), .B2(n26726), .A1(n26705), .O(n14858) );
  MUX2S U20230 ( .A(n28534), .B(n26724), .S(gray_img[219]), .O(n26705) );
  AO12S U20231 ( .B1(n15927), .B2(n26841), .A1(n26718), .O(n14859) );
  AO12S U20232 ( .B1(n15927), .B2(n26883), .A1(n26875), .O(n14860) );
  MUX2S U20233 ( .A(n28534), .B(n26881), .S(gray_img[203]), .O(n26875) );
  ND2S U20234 ( .I1(n19897), .I2(n19896), .O(n14861) );
  MUX2S U20235 ( .A(n30056), .B(n20631), .S(gray_img[195]), .O(n19896) );
  MUX2S U20236 ( .A(n29597), .B(n20082), .S(gray_img[123]), .O(n19522) );
  ND2S U20237 ( .I1(n19751), .I2(n19750), .O(n14863) );
  ND2S U20238 ( .I1(n15880), .I2(n20499), .O(n19751) );
  MUX2S U20239 ( .A(n30056), .B(n20499), .S(gray_img[115]), .O(n19750) );
  MUX2S U20240 ( .A(n29597), .B(n20617), .S(gray_img[107]), .O(n19855) );
  AO12S U20241 ( .B1(n15927), .B2(n27545), .A1(n27386), .O(n14865) );
  MUX2S U20242 ( .A(n15889), .B(n27543), .S(gray_img[99]), .O(n27386) );
  AO12S U20243 ( .B1(n15927), .B2(n26709), .A1(n26700), .O(n14866) );
  MUX2S U20244 ( .A(n28534), .B(n26707), .S(gray_img[91]), .O(n26700) );
  AO12S U20245 ( .B1(n15927), .B2(n26722), .A1(n26713), .O(n14867) );
  MUX2S U20246 ( .A(n28534), .B(n26720), .S(gray_img[83]), .O(n26713) );
  AO12S U20247 ( .B1(n15880), .B2(n26879), .A1(n26870), .O(n14868) );
  MUX2S U20248 ( .A(n27447), .B(n26877), .S(gray_img[75]), .O(n26870) );
  ND2S U20249 ( .I1(n20630), .I2(n20629), .O(n14869) );
  ND2S U20250 ( .I1(n15880), .I2(n20628), .O(n20630) );
  ND2S U20251 ( .I1(n21560), .I2(n21559), .O(n15812) );
  ND2S U20252 ( .I1(n30120), .I2(n23458), .O(n23461) );
  AO12S U20253 ( .B1(n28847), .B2(n28790), .A1(n28789), .O(n14875) );
  ND2S U20254 ( .I1(n28530), .I2(n28840), .O(n28786) );
  MUX2S U20255 ( .A(n30044), .B(n28840), .S(gray_img[140]), .O(n28787) );
  ND2S U20256 ( .I1(n28727), .I2(n28221), .O(n28224) );
  OA12S U20257 ( .B1(n29837), .B2(n28730), .A1(n28222), .O(n28223) );
  MUX2S U20258 ( .A(n15904), .B(n28728), .S(gray_img[412]), .O(n28222) );
  AO12S U20259 ( .B1(n28724), .B2(n26062), .A1(n26061), .O(n13625) );
  ND2S U20260 ( .I1(n28530), .I2(n28718), .O(n26058) );
  MUX2S U20261 ( .A(n15904), .B(n28718), .S(gray_img[956]), .O(n26059) );
  AO12S U20262 ( .B1(n26096), .B2(n25917), .A1(n25916), .O(n13626) );
  ND2S U20263 ( .I1(n28530), .I2(n26090), .O(n25913) );
  MUX2S U20264 ( .A(n15904), .B(n26090), .S(gray_img[948]), .O(n25914) );
  ND2S U20265 ( .I1(n28806), .I2(n28690), .O(n28693) );
  MUX2S U20266 ( .A(n30056), .B(n28807), .S(gray_img[404]), .O(n28691) );
  AO12S U20267 ( .B1(n25619), .B2(n25592), .A1(n25591), .O(n13627) );
  ND2S U20268 ( .I1(n28530), .I2(n25612), .O(n25588) );
  MUX2S U20269 ( .A(n29587), .B(n25612), .S(gray_img[940]), .O(n25589) );
  AO12S U20270 ( .B1(n25758), .B2(n25729), .A1(n25728), .O(n13628) );
  MUX2S U20271 ( .A(n29566), .B(n25751), .S(gray_img[932]), .O(n25726) );
  ND2S U20272 ( .I1(n28530), .I2(n25751), .O(n25725) );
  AO12S U20273 ( .B1(n30128), .B2(n30049), .A1(n30048), .O(n15069) );
  ND2S U20274 ( .I1(n28530), .I2(n30121), .O(n30045) );
  MUX2S U20275 ( .A(n30044), .B(n30121), .S(gray_img[132]), .O(n30046) );
  AO12S U20276 ( .B1(n30038), .B2(n29363), .A1(n29362), .O(n14874) );
  ND2S U20277 ( .I1(n28530), .I2(n30032), .O(n29359) );
  MUX2S U20278 ( .A(n30050), .B(n30032), .S(gray_img[396]), .O(n29360) );
  ND2S U20279 ( .I1(n30020), .I2(n29167), .O(n29170) );
  OA12S U20280 ( .B1(n29837), .B2(n30023), .A1(n29168), .O(n29169) );
  MUX2S U20281 ( .A(n30056), .B(n30021), .S(gray_img[916]), .O(n29168) );
  AO12S U20282 ( .B1(n30109), .B2(n29980), .A1(n29979), .O(n13634) );
  ND2S U20283 ( .I1(n28530), .I2(n30103), .O(n29976) );
  MUX2S U20284 ( .A(n29597), .B(n30103), .S(gray_img[388]), .O(n29977) );
  ND2S U20285 ( .I1(n28247), .I2(n28186), .O(n28189) );
  OA12S U20286 ( .B1(n29837), .B2(n28250), .A1(n28187), .O(n28188) );
  MUX2S U20287 ( .A(n30005), .B(n28248), .S(gray_img[284]), .O(n28187) );
  OA12S U20288 ( .B1(n29837), .B2(n28709), .A1(n28655), .O(n28656) );
  MUX2S U20289 ( .A(n15904), .B(n28707), .S(gray_img[276]), .O(n28655) );
  AO12S U20290 ( .B1(n29381), .B2(n29329), .A1(n29328), .O(n13703) );
  ND2S U20291 ( .I1(n28530), .I2(n29374), .O(n29325) );
  MUX2S U20292 ( .A(n29597), .B(n29374), .S(gray_img[268]), .O(n29326) );
  AO12S U20293 ( .B1(n30012), .B2(n29955), .A1(n29954), .O(n13732) );
  ND2S U20294 ( .I1(n28530), .I2(n30006), .O(n29951) );
  MUX2S U20295 ( .A(n30005), .B(n30006), .S(gray_img[260]), .O(n29952) );
  AO12S U20296 ( .B1(n30087), .B2(n28829), .A1(n28828), .O(n13750) );
  ND2S U20297 ( .I1(n28530), .I2(n30081), .O(n28825) );
  MUX2S U20298 ( .A(n15904), .B(n30081), .S(gray_img[12]), .O(n28826) );
  AO12S U20299 ( .B1(n27851), .B2(n27803), .A1(n27802), .O(n13758) );
  ND2S U20300 ( .I1(n28530), .I2(n27845), .O(n27799) );
  MUX2S U20301 ( .A(n29566), .B(n27845), .S(gray_img[156]), .O(n27800) );
  AO12S U20302 ( .B1(n30076), .B2(n27313), .A1(n27312), .O(n13768) );
  ND2S U20303 ( .I1(n28530), .I2(n30070), .O(n27309) );
  MUX2S U20304 ( .A(n30056), .B(n30070), .S(gray_img[148]), .O(n27310) );
  AO12S U20305 ( .B1(n27821), .B2(n27761), .A1(n27760), .O(n13788) );
  ND2S U20306 ( .I1(n28530), .I2(n27814), .O(n27757) );
  MUX2S U20307 ( .A(n30005), .B(n27814), .S(gray_img[28]), .O(n27758) );
  AO12S U20308 ( .B1(n27378), .B2(n27339), .A1(n27338), .O(n13798) );
  ND2S U20309 ( .I1(n28530), .I2(n27371), .O(n27335) );
  AO12S U20310 ( .B1(n30098), .B2(n29466), .A1(n29465), .O(n13841) );
  ND2S U20311 ( .I1(n28530), .I2(n30092), .O(n29462) );
  MUX2S U20312 ( .A(n29566), .B(n30092), .S(gray_img[900]), .O(n29463) );
  AO12S U20313 ( .B1(n26080), .B2(n26034), .A1(n26033), .O(n13863) );
  ND2S U20314 ( .I1(n28530), .I2(n26073), .O(n26030) );
  MUX2S U20315 ( .A(n15904), .B(n26073), .S(gray_img[828]), .O(n26031) );
  AO12S U20316 ( .B1(n25936), .B2(n25886), .A1(n25885), .O(n13869) );
  ND2S U20317 ( .I1(n28530), .I2(n25929), .O(n25882) );
  MUX2S U20318 ( .A(n25928), .B(n25929), .S(gray_img[820]), .O(n25883) );
  AO12S U20319 ( .B1(n25750), .B2(n25704), .A1(n25703), .O(n13881) );
  ND2S U20320 ( .I1(n28530), .I2(n25744), .O(n25700) );
  MUX2S U20321 ( .A(n25928), .B(n25744), .S(gray_img[804]), .O(n25701) );
  AO12S U20322 ( .B1(n29273), .B2(n29247), .A1(n29246), .O(n13887) );
  ND2S U20323 ( .I1(n28530), .I2(n29266), .O(n29243) );
  MUX2S U20324 ( .A(n30050), .B(n29266), .S(gray_img[796]), .O(n29244) );
  AO12S U20325 ( .B1(n29192), .B2(n29146), .A1(n29145), .O(n13893) );
  ND2S U20326 ( .I1(n28530), .I2(n29186), .O(n29142) );
  MUX2S U20327 ( .A(n15904), .B(n29186), .S(gray_img[788]), .O(n29143) );
  AO12S U20328 ( .B1(n29487), .B2(n29441), .A1(n29440), .O(n13905) );
  ND2S U20329 ( .I1(n28530), .I2(n29481), .O(n29437) );
  MUX2S U20330 ( .A(n30050), .B(n29481), .S(gray_img[772]), .O(n29438) );
  ND2S U20331 ( .I1(n28136), .I2(n27939), .O(n27942) );
  OA12S U20332 ( .B1(n29837), .B2(n28139), .A1(n27940), .O(n27941) );
  MUX2S U20333 ( .A(n30005), .B(n28137), .S(gray_img[700]), .O(n27940) );
  AO12S U20334 ( .B1(n28214), .B2(n28110), .A1(n28109), .O(n13933) );
  ND2S U20335 ( .I1(n28530), .I2(n28208), .O(n28106) );
  MUX2S U20336 ( .A(n30005), .B(n28208), .S(gray_img[692]), .O(n28107) );
  AO12S U20337 ( .B1(n28607), .B2(n28441), .A1(n28440), .O(n13940) );
  ND2S U20338 ( .I1(n28530), .I2(n28601), .O(n28437) );
  MUX2S U20339 ( .A(n15904), .B(n28601), .S(gray_img[684]), .O(n28438) );
  AO12S U20340 ( .B1(n28588), .B2(n28547), .A1(n28546), .O(n13947) );
  ND2S U20341 ( .I1(n28530), .I2(n28581), .O(n28543) );
  MUX2S U20342 ( .A(n30056), .B(n28581), .S(gray_img[676]), .O(n28544) );
  OA112S U20343 ( .C1(n29340), .C2(n23205), .A1(n23204), .B1(n23203), .O(
        n23206) );
  AO12S U20344 ( .B1(n29040), .B2(n28998), .A1(n28997), .O(n13963) );
  ND2S U20345 ( .I1(n28530), .I2(n29033), .O(n28994) );
  MUX2S U20346 ( .A(n29587), .B(n29033), .S(gray_img[660]), .O(n28995) );
  AO12S U20347 ( .B1(n29904), .B2(n29868), .A1(n29867), .O(n13972) );
  ND2S U20348 ( .I1(n28530), .I2(n29898), .O(n29864) );
  MUX2S U20349 ( .A(n15904), .B(n29898), .S(gray_img[652]), .O(n29865) );
  ND2S U20350 ( .I1(n29993), .I2(n29691), .O(n29694) );
  OA12S U20351 ( .B1(n29837), .B2(n29996), .A1(n29692), .O(n29693) );
  MUX2S U20352 ( .A(n15904), .B(n29994), .S(gray_img[644]), .O(n29692) );
  ND2S U20353 ( .I1(n23492), .I2(n23355), .O(n23358) );
  MUX2S U20354 ( .A(n30056), .B(n23493), .S(gray_img[572]), .O(n23356) );
  AO12S U20355 ( .B1(n28128), .B2(n28079), .A1(n28078), .O(n14015) );
  ND2S U20356 ( .I1(n28530), .I2(n28121), .O(n28075) );
  MUX2S U20357 ( .A(n30044), .B(n28121), .S(gray_img[564]), .O(n28076) );
  AO12S U20358 ( .B1(n28459), .B2(n28410), .A1(n28409), .O(n14024) );
  ND2S U20359 ( .I1(n28530), .I2(n28452), .O(n28406) );
  MUX2S U20360 ( .A(n29032), .B(n28452), .S(gray_img[556]), .O(n28407) );
  ND2S U20361 ( .I1(n28671), .I2(n28566), .O(n28569) );
  OA12S U20362 ( .B1(n29837), .B2(n28674), .A1(n28567), .O(n28568) );
  MUX2S U20363 ( .A(n15904), .B(n28672), .S(gray_img[548]), .O(n28567) );
  AO12S U20364 ( .B1(n28950), .B2(n28924), .A1(n28923), .O(n14042) );
  ND2S U20365 ( .I1(n28530), .I2(n28943), .O(n28920) );
  MUX2S U20366 ( .A(n30056), .B(n28943), .S(gray_img[540]), .O(n28921) );
  ND2S U20367 ( .I1(n29043), .I2(n29022), .O(n29025) );
  MUX2S U20368 ( .A(n30044), .B(n29044), .S(gray_img[532]), .O(n29023) );
  OA12S U20369 ( .B1(n29837), .B2(n29883), .A1(n29836), .O(n29838) );
  MUX2S U20370 ( .A(n30005), .B(n29881), .S(gray_img[524]), .O(n29836) );
  AO12S U20371 ( .B1(n26473), .B2(n26426), .A1(n26425), .O(n14094) );
  ND2S U20372 ( .I1(n28530), .I2(n26466), .O(n26422) );
  MUX2S U20373 ( .A(n15904), .B(n26466), .S(gray_img[444]), .O(n26423) );
  AO12S U20374 ( .B1(n27840), .B2(n26281), .A1(n26280), .O(n14103) );
  ND2S U20375 ( .I1(n28530), .I2(n27834), .O(n26277) );
  MUX2S U20376 ( .A(n29587), .B(n27834), .S(gray_img[436]), .O(n26278) );
  ND2S U20377 ( .I1(n23121), .I2(n23105), .O(n23108) );
  MUX2S U20378 ( .A(n29587), .B(n25151), .S(gray_img[428]), .O(n23106) );
  OA12S U20379 ( .B1(n29837), .B2(n27224), .A1(n27197), .O(n27200) );
  ND2S U20380 ( .I1(n27226), .I2(n27198), .O(n27199) );
  MUX2S U20381 ( .A(n30050), .B(n27222), .S(gray_img[420]), .O(n27197) );
  AO12S U20382 ( .B1(n26489), .B2(n26455), .A1(n26454), .O(n14138) );
  ND2S U20383 ( .I1(n28530), .I2(n26483), .O(n26451) );
  MUX2S U20384 ( .A(n29597), .B(n26483), .S(gray_img[316]), .O(n26452) );
  ND2S U20385 ( .I1(n26327), .I2(n26303), .O(n26304) );
  OA12S U20386 ( .B1(n29837), .B2(n26324), .A1(n26302), .O(n26305) );
  MUX2S U20387 ( .A(n15904), .B(n26322), .S(gray_img[308]), .O(n26302) );
  AO12S U20388 ( .B1(n27121), .B2(n27092), .A1(n27091), .O(n14156) );
  MUX2S U20389 ( .A(n29597), .B(n27114), .S(gray_img[300]), .O(n27089) );
  ND2S U20390 ( .I1(n28530), .I2(n27114), .O(n27088) );
  OA12S U20391 ( .B1(n29837), .B2(n27254), .A1(n27208), .O(n27209) );
  ND2S U20392 ( .I1(n27251), .I2(n27207), .O(n27210) );
  MUX2S U20393 ( .A(n30056), .B(n27252), .S(gray_img[292]), .O(n27208) );
  AO12S U20394 ( .B1(n27692), .B2(n27646), .A1(n27645), .O(n14182) );
  ND2S U20395 ( .I1(n28530), .I2(n27685), .O(n27642) );
  MUX2S U20396 ( .A(n30056), .B(n27685), .S(gray_img[188]), .O(n27643) );
  AO12S U20397 ( .B1(n27785), .B2(n27501), .A1(n27500), .O(n14191) );
  ND2S U20398 ( .I1(n28530), .I2(n27779), .O(n27497) );
  MUX2S U20399 ( .A(n30044), .B(n27779), .S(gray_img[180]), .O(n27498) );
  OA12S U20400 ( .B1(n29837), .B2(n27358), .A1(n26809), .O(n26810) );
  MUX2S U20401 ( .A(n30056), .B(n27356), .S(gray_img[172]), .O(n26809) );
  AO12S U20402 ( .B1(n26939), .B2(n26913), .A1(n26912), .O(n14209) );
  MUX2S U20403 ( .A(n29032), .B(n26932), .S(gray_img[164]), .O(n26910) );
  ND2S U20404 ( .I1(n28530), .I2(n26932), .O(n26909) );
  AO12S U20405 ( .B1(n27708), .B2(n27674), .A1(n27673), .O(n14226) );
  ND2S U20406 ( .I1(n28530), .I2(n27702), .O(n27670) );
  MUX2S U20407 ( .A(n30056), .B(n27702), .S(gray_img[60]), .O(n27671) );
  AO12S U20408 ( .B1(n27556), .B2(n27527), .A1(n27526), .O(n14235) );
  MUX2S U20409 ( .A(n29032), .B(n27550), .S(gray_img[52]), .O(n27524) );
  ND2S U20410 ( .I1(n28530), .I2(n27550), .O(n27523) );
  AO12S U20411 ( .B1(n26931), .B2(n26893), .A1(n26892), .O(n14253) );
  ND2S U20412 ( .I1(n28530), .I2(n26924), .O(n26889) );
  MUX2S U20413 ( .A(n29597), .B(n26924), .S(gray_img[36]), .O(n26890) );
  AO12S U20414 ( .B1(n29604), .B2(n29565), .A1(n29564), .O(n14871) );
  MUX2S U20415 ( .A(n29566), .B(n29598), .S(gray_img[908]), .O(n29562) );
  ND2S U20416 ( .I1(n28530), .I2(n29598), .O(n29561) );
  ND2S U20417 ( .I1(n28530), .I2(n20614), .O(n19410) );
  ND2S U20418 ( .I1(n28530), .I2(n20608), .O(n19795) );
  AO12S U20419 ( .B1(n28530), .B2(n25836), .A1(n25827), .O(n14880) );
  MUX2S U20420 ( .A(n27447), .B(n25834), .S(gray_img[2020]), .O(n25827) );
  AO12S U20421 ( .B1(n28530), .B2(n25473), .A1(n25463), .O(n14881) );
  MUX2S U20422 ( .A(n15889), .B(n25471), .S(gray_img[2012]), .O(n25463) );
  AO12S U20423 ( .B1(n28530), .B2(n25761), .A1(n25451), .O(n14882) );
  AO12S U20424 ( .B1(n28530), .B2(n28803), .A1(n25626), .O(n14883) );
  MUX2S U20425 ( .A(n27447), .B(n28801), .S(gray_img[1996]), .O(n25626) );
  ND2S U20426 ( .I1(n19264), .I2(n19263), .O(n14884) );
  ND2S U20427 ( .I1(n28530), .I2(n20209), .O(n19263) );
  ND2S U20428 ( .I1(n28530), .I2(n20746), .O(n19352) );
  MUX2S U20429 ( .A(n29566), .B(n20746), .S(gray_img[1980]), .O(n19351) );
  ND2S U20430 ( .I1(n28530), .I2(n20849), .O(n19393) );
  MUX2S U20431 ( .A(n29597), .B(n20849), .S(gray_img[1972]), .O(n19394) );
  ND2S U20432 ( .I1(n19270), .I2(n19269), .O(n14887) );
  ND2S U20433 ( .I1(n28530), .I2(n20202), .O(n19269) );
  ND2S U20434 ( .I1(n20327), .I2(n20326), .O(n14888) );
  ND2S U20435 ( .I1(n28530), .I2(n20586), .O(n20326) );
  ND2S U20436 ( .I1(n19286), .I2(n19285), .O(n14889) );
  MUX2S U20437 ( .A(n29566), .B(n19970), .S(gray_img[1948]), .O(n19286) );
  ND2S U20438 ( .I1(n28530), .I2(n19970), .O(n19285) );
  ND2S U20439 ( .I1(n19304), .I2(n19303), .O(n14890) );
  ND2S U20440 ( .I1(n28530), .I2(n20389), .O(n19303) );
  MUX2S U20441 ( .A(n30056), .B(n20389), .S(gray_img[1940]), .O(n19304) );
  ND2S U20442 ( .I1(n28530), .I2(n20424), .O(n19230) );
  MUX2S U20443 ( .A(n30044), .B(n20424), .S(gray_img[1932]), .O(n19229) );
  ND2S U20444 ( .I1(n19300), .I2(n19299), .O(n14892) );
  ND2S U20445 ( .I1(n28530), .I2(n20373), .O(n19299) );
  MUX2S U20446 ( .A(n20842), .B(n20373), .S(gray_img[1924]), .O(n19300) );
  ND2S U20447 ( .I1(n28530), .I2(n20430), .O(n19228) );
  MUX2S U20448 ( .A(n30056), .B(n20430), .S(gray_img[1916]), .O(n19227) );
  ND2S U20449 ( .I1(n28530), .I2(n20063), .O(n19248) );
  ND2S U20450 ( .I1(n28530), .I2(n20544), .O(n19218) );
  MUX2S U20451 ( .A(n30044), .B(n20544), .S(gray_img[1900]), .O(n19217) );
  AO12S U20452 ( .B1(n28530), .B2(n25832), .A1(n25822), .O(n14896) );
  MUX2S U20453 ( .A(n27447), .B(n25830), .S(gray_img[1892]), .O(n25822) );
  AO12S U20454 ( .B1(n28530), .B2(n25477), .A1(n25468), .O(n14897) );
  AO12S U20455 ( .B1(n28530), .B2(n25460), .A1(n25455), .O(n14898) );
  AO12S U20456 ( .B1(n28530), .B2(n25631), .A1(n25621), .O(n14899) );
  MUX2S U20457 ( .A(n15889), .B(n25629), .S(gray_img[1868]), .O(n25621) );
  MUX2S U20458 ( .A(n29566), .B(n20504), .S(gray_img[1860]), .O(n19215) );
  ND2S U20459 ( .I1(n28530), .I2(n20504), .O(n19216) );
  ND2S U20460 ( .I1(n28530), .I2(n20740), .O(n19368) );
  MUX2S U20461 ( .A(n29566), .B(n20740), .S(gray_img[1852]), .O(n19367) );
  ND2S U20462 ( .I1(n28530), .I2(n20862), .O(n19377) );
  MUX2S U20463 ( .A(n29597), .B(n20862), .S(gray_img[1844]), .O(n19378) );
  ND2S U20464 ( .I1(n19268), .I2(n19267), .O(n14903) );
  ND2S U20465 ( .I1(n28530), .I2(n20142), .O(n19267) );
  ND2S U20466 ( .I1(n19276), .I2(n19275), .O(n14904) );
  ND2S U20467 ( .I1(n28530), .I2(n20156), .O(n19275) );
  ND2S U20468 ( .I1(n19282), .I2(n19281), .O(n14905) );
  ND2S U20469 ( .I1(n28530), .I2(n20296), .O(n19281) );
  MUX2S U20470 ( .A(n29587), .B(n20296), .S(gray_img[1820]), .O(n19282) );
  ND2S U20471 ( .I1(n20339), .I2(n20338), .O(n14906) );
  ND2S U20472 ( .I1(n28530), .I2(n20354), .O(n20338) );
  MUX2S U20473 ( .A(n29566), .B(n20354), .S(gray_img[1812]), .O(n20339) );
  ND2S U20474 ( .I1(n28530), .I2(n20319), .O(n19206) );
  MUX2S U20475 ( .A(n30044), .B(n20319), .S(gray_img[1804]), .O(n19205) );
  ND2S U20476 ( .I1(n19310), .I2(n19309), .O(n14908) );
  MUX2S U20477 ( .A(n29597), .B(n20376), .S(gray_img[1796]), .O(n19310) );
  ND2S U20478 ( .I1(n28530), .I2(n20376), .O(n19309) );
  MUX2S U20479 ( .A(n29566), .B(n20547), .S(gray_img[1788]), .O(n19231) );
  ND2S U20480 ( .I1(n28530), .I2(n20547), .O(n19232) );
  MUX2S U20481 ( .A(n29566), .B(n20541), .S(gray_img[1780]), .O(n19237) );
  ND2S U20482 ( .I1(n28530), .I2(n20541), .O(n19238) );
  ND2S U20483 ( .I1(n28530), .I2(n20449), .O(n19246) );
  MUX2S U20484 ( .A(n30050), .B(n20449), .S(gray_img[1772]), .O(n19245) );
  AO12S U20485 ( .B1(n28530), .B2(n25778), .A1(n25768), .O(n14912) );
  AO12S U20486 ( .B1(n28530), .B2(n25510), .A1(n25500), .O(n14913) );
  AO12S U20487 ( .B1(n28530), .B2(n25498), .A1(n25489), .O(n14914) );
  MUX2S U20488 ( .A(n15889), .B(n25496), .S(gray_img[1748]), .O(n25489) );
  AO12S U20489 ( .B1(n28530), .B2(n25649), .A1(n25639), .O(n14915) );
  MUX2S U20490 ( .A(n27447), .B(n25647), .S(gray_img[1740]), .O(n25639) );
  MUX2S U20491 ( .A(n29597), .B(n19955), .S(gray_img[1732]), .O(n19233) );
  ND2S U20492 ( .I1(n28530), .I2(n19955), .O(n19234) );
  ND2S U20493 ( .I1(n28530), .I2(n20737), .O(n19356) );
  MUX2S U20494 ( .A(n30044), .B(n20737), .S(gray_img[1724]), .O(n19355) );
  ND2S U20495 ( .I1(n28530), .I2(n20846), .O(n19371) );
  MUX2S U20496 ( .A(n20830), .B(n20846), .S(gray_img[1716]), .O(n19372) );
  ND2S U20497 ( .I1(n28530), .I2(n20827), .O(n19389) );
  MUX2S U20498 ( .A(n30050), .B(n20827), .S(gray_img[1708]), .O(n19390) );
  ND2S U20499 ( .I1(n28530), .I2(n20787), .O(n19379) );
  MUX2S U20500 ( .A(n30056), .B(n20787), .S(gray_img[1700]), .O(n19380) );
  ND2S U20501 ( .I1(n19256), .I2(n19255), .O(n14921) );
  ND2S U20502 ( .I1(n28530), .I2(n20599), .O(n19255) );
  MUX2S U20503 ( .A(n30044), .B(n20599), .S(gray_img[1692]), .O(n19256) );
  ND2S U20504 ( .I1(n19266), .I2(n19265), .O(n14922) );
  ND2S U20505 ( .I1(n28530), .I2(n20605), .O(n19265) );
  MUX2S U20506 ( .A(n30044), .B(n20605), .S(gray_img[1684]), .O(n19266) );
  ND2S U20507 ( .I1(n28530), .I2(n20531), .O(n19210) );
  MUX2S U20508 ( .A(n29566), .B(n20531), .S(gray_img[1676]), .O(n19209) );
  ND2S U20509 ( .I1(n19254), .I2(n19253), .O(n14924) );
  ND2S U20510 ( .I1(n28530), .I2(n20583), .O(n19253) );
  MUX2S U20511 ( .A(n29597), .B(n20583), .S(gray_img[1668]), .O(n19254) );
  ND2S U20512 ( .I1(n28530), .I2(n20509), .O(n19226) );
  MUX2S U20513 ( .A(n29597), .B(n20525), .S(gray_img[1652]), .O(n19213) );
  ND2S U20514 ( .I1(n28530), .I2(n20525), .O(n19214) );
  ND2S U20515 ( .I1(n28530), .I2(n20463), .O(n19222) );
  AO12S U20516 ( .B1(n28530), .B2(n25899), .A1(n25773), .O(n14928) );
  MUX2S U20517 ( .A(n27447), .B(n25897), .S(gray_img[1636]), .O(n25773) );
  AO12S U20518 ( .B1(n28530), .B2(n25576), .A1(n25505), .O(n14929) );
  AO12S U20519 ( .B1(n28530), .B2(n25494), .A1(n25484), .O(n14930) );
  AO12S U20520 ( .B1(n28530), .B2(n25653), .A1(n25644), .O(n14931) );
  MUX2S U20521 ( .A(n29597), .B(n20528), .S(gray_img[1604]), .O(n19219) );
  ND2S U20522 ( .I1(n28530), .I2(n20528), .O(n19220) );
  ND2S U20523 ( .I1(n28530), .I2(n20731), .O(n19358) );
  MUX2S U20524 ( .A(n30056), .B(n20731), .S(gray_img[1596]), .O(n19357) );
  ND2S U20525 ( .I1(n28530), .I2(n20839), .O(n19387) );
  MUX2S U20526 ( .A(n20830), .B(n20839), .S(gray_img[1588]), .O(n19388) );
  ND2S U20527 ( .I1(n28530), .I2(n20395), .O(n19373) );
  MUX2S U20528 ( .A(n30050), .B(n20395), .S(gray_img[1580]), .O(n19374) );
  ND2S U20529 ( .I1(n28530), .I2(n20824), .O(n19383) );
  MUX2S U20530 ( .A(n30056), .B(n20824), .S(gray_img[1572]), .O(n19384) );
  ND2S U20531 ( .I1(n19280), .I2(n19279), .O(n14937) );
  MUX2S U20532 ( .A(n29587), .B(n20596), .S(gray_img[1564]), .O(n19280) );
  ND2S U20533 ( .I1(n28530), .I2(n20596), .O(n19279) );
  ND2S U20534 ( .I1(n19252), .I2(n19251), .O(n14938) );
  ND2S U20535 ( .I1(n28530), .I2(n20602), .O(n19251) );
  MUX2S U20536 ( .A(n29566), .B(n20602), .S(gray_img[1556]), .O(n19252) );
  ND2S U20537 ( .I1(n28530), .I2(n20550), .O(n19212) );
  ND2S U20538 ( .I1(n20874), .I2(n20873), .O(n14940) );
  MUX2S U20539 ( .A(n29587), .B(n20881), .S(gray_img[1540]), .O(n20874) );
  ND2S U20540 ( .I1(n28530), .I2(n20881), .O(n20873) );
  ND2S U20541 ( .I1(n28530), .I2(n20556), .O(n19204) );
  MUX2S U20542 ( .A(n30044), .B(n20556), .S(gray_img[1532]), .O(n19203) );
  ND2S U20543 ( .I1(n19182), .I2(n19181), .O(n14942) );
  ND2S U20544 ( .I1(n28530), .I2(n20512), .O(n19182) );
  ND2S U20545 ( .I1(n28530), .I2(n20440), .O(n19370) );
  MUX2S U20546 ( .A(n30050), .B(n20440), .S(gray_img[1516]), .O(n19369) );
  AO12S U20547 ( .B1(n28530), .B2(n27971), .A1(n27966), .O(n14944) );
  MUX2S U20548 ( .A(n28534), .B(n27969), .S(gray_img[1508]), .O(n27966) );
  AO12S U20549 ( .B1(n28530), .B2(n28355), .A1(n28345), .O(n14945) );
  AO12S U20550 ( .B1(n28530), .B2(n28342), .A1(n28332), .O(n14946) );
  MUX2S U20551 ( .A(n28534), .B(n28340), .S(gray_img[1492]), .O(n28332) );
  AO12S U20552 ( .B1(n28530), .B2(n28560), .A1(n28529), .O(n14947) );
  ND2S U20553 ( .I1(n28530), .I2(n20684), .O(n19348) );
  MUX2S U20554 ( .A(n30056), .B(n20684), .S(gray_img[1476]), .O(n19347) );
  ND2S U20555 ( .I1(n19978), .I2(n19977), .O(n14949) );
  ND2S U20556 ( .I1(n28530), .I2(n20709), .O(n19978) );
  ND2S U20557 ( .I1(n28530), .I2(n20821), .O(n19987) );
  MUX2S U20558 ( .A(n30044), .B(n20821), .S(gray_img[1460]), .O(n19988) );
  ND2S U20559 ( .I1(n28530), .I2(n20814), .O(n19381) );
  MUX2S U20560 ( .A(n29566), .B(n20814), .S(gray_img[1452]), .O(n19382) );
  ND2S U20561 ( .I1(n28530), .I2(n20811), .O(n19375) );
  ND2S U20562 ( .I1(n19290), .I2(n19289), .O(n14953) );
  ND2S U20563 ( .I1(n28530), .I2(n20293), .O(n19289) );
  MUX2S U20564 ( .A(n30050), .B(n20293), .S(gray_img[1436]), .O(n19290) );
  ND2S U20565 ( .I1(n19260), .I2(n19259), .O(n14954) );
  ND2S U20566 ( .I1(n28530), .I2(n20193), .O(n19259) );
  MUX2S U20567 ( .A(n20842), .B(n20193), .S(gray_img[1428]), .O(n19260) );
  ND2S U20568 ( .I1(n19194), .I2(n19193), .O(n14955) );
  ND2S U20569 ( .I1(n28530), .I2(n20035), .O(n19194) );
  ND2S U20570 ( .I1(n19278), .I2(n19277), .O(n14956) );
  ND2S U20571 ( .I1(n28530), .I2(n20359), .O(n19277) );
  MUX2S U20572 ( .A(n20842), .B(n20359), .S(gray_img[1412]), .O(n19278) );
  ND2S U20573 ( .I1(n28530), .I2(n20571), .O(n19184) );
  MUX2S U20574 ( .A(n30050), .B(n20571), .S(gray_img[1404]), .O(n19183) );
  ND2S U20575 ( .I1(n19192), .I2(n19191), .O(n14958) );
  ND2S U20576 ( .I1(n28530), .I2(n20517), .O(n19192) );
  ND2S U20577 ( .I1(n28530), .I2(n20722), .O(n19354) );
  MUX2S U20578 ( .A(n30050), .B(n20722), .S(gray_img[1388]), .O(n19353) );
  AO12S U20579 ( .B1(n28530), .B2(n28203), .A1(n27962), .O(n14960) );
  MUX2S U20580 ( .A(n28534), .B(n28201), .S(gray_img[1380]), .O(n27962) );
  AO12S U20581 ( .B1(n28530), .B2(n28359), .A1(n28350), .O(n14961) );
  MUX2S U20582 ( .A(n28534), .B(n28357), .S(gray_img[1372]), .O(n28350) );
  AO12S U20583 ( .B1(n28530), .B2(n28596), .A1(n28337), .O(n14962) );
  MUX2S U20584 ( .A(n15889), .B(n28594), .S(gray_img[1364]), .O(n28337) );
  AO12S U20585 ( .B1(n28530), .B2(n28536), .A1(n28524), .O(n14963) );
  ND2S U20586 ( .I1(n28530), .I2(n20734), .O(n19982) );
  MUX2S U20587 ( .A(n30044), .B(n20734), .S(gray_img[1348]), .O(n19981) );
  ND2S U20588 ( .I1(n28530), .I2(n20695), .O(n19976) );
  MUX2S U20589 ( .A(n30050), .B(n20695), .S(gray_img[1340]), .O(n19975) );
  ND2S U20590 ( .I1(n28530), .I2(n20833), .O(n19989) );
  MUX2S U20591 ( .A(n30056), .B(n20833), .S(gray_img[1332]), .O(n19990) );
  ND2S U20592 ( .I1(n28530), .I2(n20836), .O(n19391) );
  MUX2S U20593 ( .A(n29566), .B(n20836), .S(gray_img[1324]), .O(n19392) );
  ND2S U20594 ( .I1(n28530), .I2(n20843), .O(n19385) );
  MUX2S U20595 ( .A(n29597), .B(n20843), .S(gray_img[1316]), .O(n19386) );
  ND2S U20596 ( .I1(n19274), .I2(n19273), .O(n14969) );
  ND2S U20597 ( .I1(n28530), .I2(n20129), .O(n19273) );
  ND2S U20598 ( .I1(n19284), .I2(n19283), .O(n14970) );
  ND2S U20599 ( .I1(n28530), .I2(n20362), .O(n19283) );
  MUX2S U20600 ( .A(n15904), .B(n20362), .S(gray_img[1300]), .O(n19284) );
  ND2S U20601 ( .I1(n19200), .I2(n19199), .O(n14971) );
  ND2S U20602 ( .I1(n28530), .I2(n20427), .O(n19200) );
  ND2S U20603 ( .I1(n19288), .I2(n19287), .O(n14972) );
  ND2S U20604 ( .I1(n28530), .I2(n20392), .O(n19287) );
  MUX2S U20605 ( .A(n30050), .B(n20392), .S(gray_img[1284]), .O(n19288) );
  ND2S U20606 ( .I1(n28530), .I2(n20655), .O(n19362) );
  MUX2S U20607 ( .A(n20808), .B(n20655), .S(gray_img[1276]), .O(n19361) );
  ND2S U20608 ( .I1(n28530), .I2(n20725), .O(n19986) );
  MUX2S U20609 ( .A(n20808), .B(n20725), .S(gray_img[1268]), .O(n19985) );
  ND2S U20610 ( .I1(n28530), .I2(n20719), .O(n19360) );
  MUX2S U20611 ( .A(n30044), .B(n20719), .S(gray_img[1260]), .O(n19359) );
  AO12S U20612 ( .B1(n28530), .B2(n28031), .A1(n28025), .O(n14976) );
  AO12S U20613 ( .B1(n28530), .B2(n28288), .A1(n28279), .O(n14977) );
  AO12S U20614 ( .B1(n28530), .B2(n28271), .A1(n28261), .O(n14978) );
  MUX2S U20615 ( .A(n28534), .B(n28269), .S(gray_img[1236]), .O(n28261) );
  AO12S U20616 ( .B1(n28530), .B2(n28475), .A1(n28466), .O(n14979) );
  ND2S U20617 ( .I1(n28530), .I2(n20702), .O(n19980) );
  MUX2S U20618 ( .A(n29587), .B(n20702), .S(gray_img[1220]), .O(n19979) );
  ND2S U20619 ( .I1(n19733), .I2(n19732), .O(n14981) );
  ND2S U20620 ( .I1(n28530), .I2(n20757), .O(n19733) );
  MUX2S U20621 ( .A(n30044), .B(n20757), .S(gray_img[1212]), .O(n19732) );
  ND2S U20622 ( .I1(n28530), .I2(n20857), .O(n19993) );
  MUX2S U20623 ( .A(n30044), .B(n20857), .S(gray_img[1204]), .O(n19994) );
  ND2S U20624 ( .I1(n28530), .I2(n20435), .O(n19669) );
  MUX2S U20625 ( .A(n29587), .B(n20435), .S(gray_img[1196]), .O(n19668) );
  ND2S U20626 ( .I1(n19292), .I2(n19291), .O(n14984) );
  MUX2S U20627 ( .A(n29566), .B(n20379), .S(gray_img[1188]), .O(n19292) );
  ND2S U20628 ( .I1(n28530), .I2(n20379), .O(n19291) );
  ND2S U20629 ( .I1(n19298), .I2(n19297), .O(n14985) );
  ND2S U20630 ( .I1(n28530), .I2(n20159), .O(n19297) );
  MUX2S U20631 ( .A(n29597), .B(n20159), .S(gray_img[1180]), .O(n19298) );
  ND2S U20632 ( .I1(n28530), .I2(n20316), .O(n19763) );
  MUX2S U20633 ( .A(n29597), .B(n20316), .S(gray_img[1172]), .O(n19762) );
  MUX2S U20634 ( .A(n29597), .B(n20553), .S(gray_img[1164]), .O(n19179) );
  ND2S U20635 ( .I1(n28530), .I2(n20553), .O(n19180) );
  ND2S U20636 ( .I1(n28530), .I2(n20240), .O(n19705) );
  MUX2S U20637 ( .A(n29566), .B(n20240), .S(gray_img[1156]), .O(n19704) );
  ND2S U20638 ( .I1(n28530), .I2(n20716), .O(n19366) );
  MUX2S U20639 ( .A(n30044), .B(n20716), .S(gray_img[1148]), .O(n19365) );
  ND2S U20640 ( .I1(n28530), .I2(n20124), .O(n19984) );
  MUX2S U20641 ( .A(n20808), .B(n20124), .S(gray_img[1140]), .O(n19983) );
  ND2S U20642 ( .I1(n28530), .I2(n20728), .O(n19364) );
  MUX2S U20643 ( .A(n30056), .B(n20728), .S(gray_img[1132]), .O(n19363) );
  AO12S U20644 ( .B1(n28530), .B2(n28092), .A1(n28020), .O(n14992) );
  MUX2S U20645 ( .A(n28534), .B(n28090), .S(gray_img[1124]), .O(n28020) );
  AO12S U20646 ( .B1(n28530), .B2(n28284), .A1(n28274), .O(n14993) );
  MUX2S U20647 ( .A(n28534), .B(n28282), .S(gray_img[1116]), .O(n28274) );
  AO12S U20648 ( .B1(n28530), .B2(n28423), .A1(n28266), .O(n14994) );
  AO12S U20649 ( .B1(n28530), .B2(n28480), .A1(n28477), .O(n14995) );
  ND2S U20650 ( .I1(n28530), .I2(n20743), .O(n19350) );
  MUX2S U20651 ( .A(n30050), .B(n20743), .S(gray_img[1092]), .O(n19349) );
  ND2S U20652 ( .I1(n19728), .I2(n19727), .O(n14997) );
  ND2S U20653 ( .I1(n28530), .I2(n20760), .O(n19728) );
  MUX2S U20654 ( .A(n30056), .B(n20760), .S(gray_img[1084]), .O(n19727) );
  ND2S U20655 ( .I1(n28530), .I2(n20854), .O(n19991) );
  MUX2S U20656 ( .A(n30044), .B(n20854), .S(gray_img[1076]), .O(n19992) );
  ND2S U20657 ( .I1(n28530), .I2(n20611), .O(n19673) );
  MUX2S U20658 ( .A(n29587), .B(n20611), .S(gray_img[1068]), .O(n19672) );
  ND2S U20659 ( .I1(n19296), .I2(n19295), .O(n15000) );
  MUX2S U20660 ( .A(n29587), .B(n20368), .S(gray_img[1060]), .O(n19296) );
  ND2S U20661 ( .I1(n28530), .I2(n20368), .O(n19295) );
  ND2S U20662 ( .I1(n19294), .I2(n19293), .O(n15001) );
  ND2S U20663 ( .I1(n28530), .I2(n20184), .O(n19293) );
  MUX2S U20664 ( .A(n29587), .B(n20184), .S(gray_img[1052]), .O(n19294) );
  ND2S U20665 ( .I1(n19775), .I2(n19774), .O(n15002) );
  ND2S U20666 ( .I1(n28530), .I2(n20255), .O(n19775) );
  MUX2S U20667 ( .A(n29587), .B(n20255), .S(gray_img[1044]), .O(n19774) );
  ND2S U20668 ( .I1(n28530), .I2(n20235), .O(n19421) );
  MUX2S U20669 ( .A(n29566), .B(n20235), .S(gray_img[1036]), .O(n19420) );
  ND2S U20670 ( .I1(n28530), .I2(n20311), .O(n19698) );
  ND2S U20671 ( .I1(n28530), .I2(n20099), .O(n19178) );
  ND2S U20672 ( .I1(n28530), .I2(n20562), .O(n19196) );
  ND2S U20673 ( .I1(n19306), .I2(n19305), .O(n15007) );
  ND2S U20674 ( .I1(n28530), .I2(n20384), .O(n19305) );
  AO12S U20675 ( .B1(n28530), .B2(n27829), .A1(n26219), .O(n15008) );
  MUX2S U20676 ( .A(n28534), .B(n27827), .S(gray_img[996]), .O(n26219) );
  AO12S U20677 ( .B1(n28530), .B2(n27081), .A1(n27071), .O(n15009) );
  AO12S U20678 ( .B1(n28530), .B2(n27065), .A1(n27055), .O(n15010) );
  MUX2S U20679 ( .A(n27447), .B(n27063), .S(gray_img[980]), .O(n27055) );
  AO12S U20680 ( .B1(n28530), .B2(n27261), .A1(n27185), .O(n15011) );
  MUX2S U20681 ( .A(n27447), .B(n27259), .S(gray_img[972]), .O(n27185) );
  ND2S U20682 ( .I1(n19258), .I2(n19257), .O(n15012) );
  ND2S U20683 ( .I1(n28530), .I2(n20580), .O(n19257) );
  MUX2S U20684 ( .A(n29587), .B(n20580), .S(gray_img[964]), .O(n19258) );
  ND2S U20685 ( .I1(n28530), .I2(n20452), .O(n19190) );
  ND2S U20686 ( .I1(n28530), .I2(n20559), .O(n19186) );
  ND2S U20687 ( .I1(n19272), .I2(n19271), .O(n15015) );
  ND2S U20688 ( .I1(n28530), .I2(n20212), .O(n19271) );
  AO12S U20689 ( .B1(n28530), .B2(n26224), .A1(n26214), .O(n15016) );
  MUX2S U20690 ( .A(n27447), .B(n26222), .S(gray_img[868]), .O(n26214) );
  AO12S U20691 ( .B1(n28530), .B2(n30065), .A1(n27076), .O(n15017) );
  AO12S U20692 ( .B1(n28530), .B2(n27069), .A1(n27060), .O(n15018) );
  AO12S U20693 ( .B1(n28530), .B2(n27190), .A1(n27181), .O(n15019) );
  MUX2S U20694 ( .A(n28534), .B(n27188), .S(gray_img[844]), .O(n27181) );
  ND2S U20695 ( .I1(n19921), .I2(n19920), .O(n15020) );
  ND2S U20696 ( .I1(n28530), .I2(n20634), .O(n19921) );
  MUX2S U20697 ( .A(n20634), .B(n20830), .S(n22984), .O(n19920) );
  ND2S U20698 ( .I1(n28530), .I2(n20568), .O(n19188) );
  ND2S U20699 ( .I1(n28530), .I2(n20054), .O(n19202) );
  ND2S U20700 ( .I1(n19262), .I2(n19261), .O(n15023) );
  ND2S U20701 ( .I1(n28530), .I2(n20365), .O(n19261) );
  AO12S U20702 ( .B1(n28530), .B2(n26155), .A1(n26146), .O(n15024) );
  MUX2S U20703 ( .A(n27447), .B(n26153), .S(gray_img[740]), .O(n26146) );
  AO12S U20704 ( .B1(n28530), .B2(n26996), .A1(n26986), .O(n15025) );
  AO12S U20705 ( .B1(n28530), .B2(n27009), .A1(n26999), .O(n15026) );
  MUX2S U20706 ( .A(n15889), .B(n27007), .S(gray_img[724]), .O(n26999) );
  AO12S U20707 ( .B1(n28530), .B2(n27243), .A1(n27128), .O(n15027) );
  ND2S U20708 ( .I1(n19871), .I2(n19870), .O(n15028) );
  MUX2S U20709 ( .A(n29032), .B(n20623), .S(gray_img[708]), .O(n19870) );
  ND2S U20710 ( .I1(n28530), .I2(n20623), .O(n19871) );
  ND2S U20711 ( .I1(n28530), .I2(n20565), .O(n19240) );
  ND2S U20712 ( .I1(n28530), .I2(n20534), .O(n19236) );
  MUX2S U20713 ( .A(n30050), .B(n20534), .S(gray_img[628]), .O(n19235) );
  ND2S U20714 ( .I1(n19835), .I2(n19834), .O(n15031) );
  ND2S U20715 ( .I1(n28530), .I2(n20274), .O(n19835) );
  MUX2S U20716 ( .A(n20274), .B(n20830), .S(n26185), .O(n19834) );
  AO12S U20717 ( .B1(n28530), .B2(n26160), .A1(n26150), .O(n15032) );
  AO12S U20718 ( .B1(n28530), .B2(n27105), .A1(n26991), .O(n15033) );
  AO12S U20719 ( .B1(n28530), .B2(n27013), .A1(n27004), .O(n15034) );
  MUX2S U20720 ( .A(n28534), .B(n27011), .S(gray_img[596]), .O(n27004) );
  AO12S U20721 ( .B1(n28530), .B2(n27133), .A1(n27123), .O(n15035) );
  MUX2S U20722 ( .A(n15889), .B(n27131), .S(gray_img[588]), .O(n27123) );
  ND2S U20723 ( .I1(n19302), .I2(n19301), .O(n15036) );
  ND2S U20724 ( .I1(n28530), .I2(n20591), .O(n19301) );
  MUX2S U20725 ( .A(n29587), .B(n20591), .S(gray_img[580]), .O(n19302) );
  ND2S U20726 ( .I1(n28530), .I2(n20472), .O(n19242) );
  MUX2S U20727 ( .A(n30050), .B(n20472), .S(gray_img[508]), .O(n19241) );
  ND2S U20728 ( .I1(n19250), .I2(n19249), .O(n15038) );
  ND2S U20729 ( .I1(n28530), .I2(n20477), .O(n19250) );
  ND2S U20730 ( .I1(n28530), .I2(n20480), .O(n19811) );
  MUX2S U20731 ( .A(n29597), .B(n20480), .S(gray_img[492]), .O(n19810) );
  AO12S U20732 ( .B1(n28530), .B2(n27774), .A1(n27443), .O(n15040) );
  MUX2S U20733 ( .A(n27447), .B(n27772), .S(gray_img[484]), .O(n27443) );
  AO12S U20734 ( .B1(n28530), .B2(n27352), .A1(n26754), .O(n15041) );
  AO12S U20735 ( .B1(n28530), .B2(n26747), .A1(n26737), .O(n15042) );
  MUX2S U20736 ( .A(n15889), .B(n26745), .S(gray_img[468]), .O(n26737) );
  AO12S U20737 ( .B1(n28530), .B2(n26942), .A1(n26856), .O(n15043) );
  ND2S U20738 ( .I1(n19878), .I2(n19877), .O(n15044) );
  ND2S U20739 ( .I1(n28530), .I2(n20483), .O(n19878) );
  ND2S U20740 ( .I1(n28530), .I2(n20486), .O(n19224) );
  ND2S U20741 ( .I1(n28530), .I2(n20522), .O(n19208) );
  ND2S U20742 ( .I1(n28530), .I2(n20491), .O(n19804) );
  MUX2S U20743 ( .A(n29566), .B(n20491), .S(gray_img[364]), .O(n19803) );
  AO12S U20744 ( .B1(n28530), .B2(n27449), .A1(n27438), .O(n15048) );
  MUX2S U20745 ( .A(n28534), .B(n27446), .S(gray_img[356]), .O(n27438) );
  AO12S U20746 ( .B1(n28530), .B2(n26759), .A1(n26749), .O(n15049) );
  MUX2S U20747 ( .A(n27447), .B(n26757), .S(gray_img[348]), .O(n26749) );
  AO12S U20748 ( .B1(n28530), .B2(n26743), .A1(n26733), .O(n15050) );
  AO12S U20749 ( .B1(n28530), .B2(n26861), .A1(n26851), .O(n15051) );
  ND2S U20750 ( .I1(n19308), .I2(n19307), .O(n15052) );
  ND2S U20751 ( .I1(n28530), .I2(n20147), .O(n19307) );
  MUX2S U20752 ( .A(n29587), .B(n20496), .S(gray_img[252]), .O(n19243) );
  ND2S U20753 ( .I1(n28530), .I2(n20496), .O(n19244) );
  ND2S U20754 ( .I1(n19718), .I2(n19717), .O(n15054) );
  ND2S U20755 ( .I1(n28530), .I2(n20260), .O(n19718) );
  MUX2S U20756 ( .A(n30050), .B(n20260), .S(gray_img[244]), .O(n19717) );
  ND2S U20757 ( .I1(n28530), .I2(n20620), .O(n19830) );
  MUX2S U20758 ( .A(n29566), .B(n20620), .S(gray_img[236]), .O(n19829) );
  AO12S U20759 ( .B1(n28530), .B2(n27390), .A1(n27380), .O(n15056) );
  MUX2S U20760 ( .A(n27447), .B(n27388), .S(gray_img[228]), .O(n27380) );
  AO12S U20761 ( .B1(n28530), .B2(n26726), .A1(n26704), .O(n15057) );
  MUX2S U20762 ( .A(n28534), .B(n26724), .S(gray_img[220]), .O(n26704) );
  AO12S U20763 ( .B1(n28530), .B2(n26841), .A1(n26717), .O(n15058) );
  AO12S U20764 ( .B1(n28530), .B2(n26883), .A1(n26874), .O(n15059) );
  ND2S U20765 ( .I1(n19895), .I2(n19894), .O(n15060) );
  ND2S U20766 ( .I1(n28530), .I2(n20631), .O(n19895) );
  MUX2S U20767 ( .A(n15904), .B(n20631), .S(gray_img[196]), .O(n19894) );
  MUX2S U20768 ( .A(n29566), .B(n20082), .S(gray_img[124]), .O(n19197) );
  ND2S U20769 ( .I1(n28530), .I2(n20082), .O(n19198) );
  ND2S U20770 ( .I1(n19723), .I2(n19722), .O(n15062) );
  ND2S U20771 ( .I1(n28530), .I2(n20499), .O(n19723) );
  MUX2S U20772 ( .A(n30044), .B(n20499), .S(gray_img[116]), .O(n19722) );
  ND2S U20773 ( .I1(n28530), .I2(n20617), .O(n19858) );
  MUX2S U20774 ( .A(n29587), .B(n20617), .S(gray_img[108]), .O(n19857) );
  AO12S U20775 ( .B1(n28530), .B2(n27545), .A1(n27385), .O(n15064) );
  MUX2S U20776 ( .A(n28534), .B(n27543), .S(gray_img[100]), .O(n27385) );
  AO12S U20777 ( .B1(n28530), .B2(n26709), .A1(n26699), .O(n15065) );
  AO12S U20778 ( .B1(n28530), .B2(n26722), .A1(n26712), .O(n15066) );
  AO12S U20779 ( .B1(n28530), .B2(n26879), .A1(n26869), .O(n15067) );
  ND2S U20780 ( .I1(n19912), .I2(n19911), .O(n15068) );
  ND2S U20781 ( .I1(n28530), .I2(n20628), .O(n19912) );
  MUX2S U20782 ( .A(n15904), .B(n20628), .S(gray_img[68]), .O(n19911) );
  ND2S U20783 ( .I1(n21775), .I2(n21774), .O(n15811) );
  ND2S U20784 ( .I1(n30120), .I2(n23452), .O(n23456) );
  AO12S U20785 ( .B1(n28847), .B2(n28785), .A1(n28784), .O(n15075) );
  ND2S U20786 ( .I1(n15891), .I2(n28840), .O(n28781) );
  MUX2S U20787 ( .A(n29566), .B(n28840), .S(gray_img[141]), .O(n28782) );
  ND2S U20788 ( .I1(n28727), .I2(n28255), .O(n28258) );
  OA12S U20789 ( .B1(n29831), .B2(n28730), .A1(n28256), .O(n28257) );
  MUX2S U20790 ( .A(n15904), .B(n28728), .S(gray_img[413]), .O(n28256) );
  AO12S U20791 ( .B1(n28724), .B2(n26057), .A1(n26056), .O(n13618) );
  MUX2S U20792 ( .A(n15904), .B(n28718), .S(gray_img[957]), .O(n26054) );
  AO12S U20793 ( .B1(n26096), .B2(n25912), .A1(n25911), .O(n13619) );
  ND2S U20794 ( .I1(n26445), .I2(n26090), .O(n25908) );
  MUX2S U20795 ( .A(n15904), .B(n26090), .S(gray_img[949]), .O(n25909) );
  ND2S U20796 ( .I1(n28806), .I2(n28685), .O(n28688) );
  MUX2S U20797 ( .A(n29597), .B(n28807), .S(gray_img[405]), .O(n28686) );
  AO12S U20798 ( .B1(n25619), .B2(n25587), .A1(n25586), .O(n13620) );
  MUX2S U20799 ( .A(n29566), .B(n25612), .S(gray_img[941]), .O(n25584) );
  AO12S U20800 ( .B1(n25758), .B2(n25724), .A1(n25723), .O(n13621) );
  ND2S U20801 ( .I1(n27751), .I2(n25751), .O(n25720) );
  MUX2S U20802 ( .A(n30050), .B(n25751), .S(gray_img[933]), .O(n25721) );
  AO12S U20803 ( .B1(n30128), .B2(n30043), .A1(n30042), .O(n13624) );
  ND2S U20804 ( .I1(n15891), .I2(n30121), .O(n30039) );
  MUX2S U20805 ( .A(n30050), .B(n30121), .S(gray_img[133]), .O(n30040) );
  AO12S U20806 ( .B1(n30109), .B2(n29975), .A1(n29974), .O(n13633) );
  ND2S U20807 ( .I1(n15891), .I2(n30103), .O(n29971) );
  MUX2S U20808 ( .A(n30044), .B(n30103), .S(gray_img[389]), .O(n29972) );
  ND2S U20809 ( .I1(n28247), .I2(n28246), .O(n28252) );
  OA12S U20810 ( .B1(n29831), .B2(n28250), .A1(n28249), .O(n28251) );
  MUX2S U20811 ( .A(n15904), .B(n28248), .S(gray_img[285]), .O(n28249) );
  OA12S U20812 ( .B1(n29831), .B2(n28709), .A1(n28650), .O(n28651) );
  MUX2S U20813 ( .A(n15904), .B(n28707), .S(gray_img[277]), .O(n28650) );
  AO12S U20814 ( .B1(n29381), .B2(n29319), .A1(n29318), .O(n13702) );
  MUX2S U20815 ( .A(n29587), .B(n29374), .S(gray_img[269]), .O(n29316) );
  AO12S U20816 ( .B1(n30012), .B2(n29950), .A1(n29949), .O(n13731) );
  ND2S U20817 ( .I1(n26828), .I2(n30006), .O(n29946) );
  MUX2S U20818 ( .A(n30005), .B(n30006), .S(gray_img[261]), .O(n29947) );
  AO12S U20819 ( .B1(n30087), .B2(n28824), .A1(n28823), .O(n13749) );
  MUX2S U20820 ( .A(n15904), .B(n30081), .S(gray_img[13]), .O(n28821) );
  AO12S U20821 ( .B1(n27851), .B2(n27798), .A1(n27797), .O(n13757) );
  AO12S U20822 ( .B1(n30076), .B2(n27308), .A1(n27307), .O(n13767) );
  MUX2S U20823 ( .A(n15904), .B(n30070), .S(gray_img[149]), .O(n27305) );
  AO12S U20824 ( .B1(n27821), .B2(n27756), .A1(n27755), .O(n13787) );
  ND2S U20825 ( .I1(n27751), .I2(n27814), .O(n27752) );
  MUX2S U20826 ( .A(n30005), .B(n27814), .S(gray_img[29]), .O(n27753) );
  AO12S U20827 ( .B1(n27378), .B2(n27334), .A1(n27333), .O(n13797) );
  MUX2S U20828 ( .A(n30005), .B(n27371), .S(gray_img[21]), .O(n27331) );
  ND2S U20829 ( .I1(n26445), .I2(n27371), .O(n27330) );
  AO12S U20830 ( .B1(n30038), .B2(n29324), .A1(n29323), .O(n15072) );
  MUX2S U20831 ( .A(n29597), .B(n30032), .S(gray_img[397]), .O(n29321) );
  ND2S U20832 ( .I1(n30020), .I2(n29162), .O(n29165) );
  OA12S U20833 ( .B1(n29831), .B2(n30023), .A1(n29163), .O(n29164) );
  MUX2S U20834 ( .A(n15904), .B(n30021), .S(gray_img[917]), .O(n29163) );
  AO12S U20835 ( .B1(n29604), .B2(n29560), .A1(n29559), .O(n13835) );
  MUX2S U20836 ( .A(n29587), .B(n29598), .S(gray_img[909]), .O(n29557) );
  ND2S U20837 ( .I1(n26445), .I2(n29598), .O(n29556) );
  AO12S U20838 ( .B1(n30098), .B2(n29461), .A1(n29460), .O(n13840) );
  MUX2S U20839 ( .A(n29597), .B(n30092), .S(gray_img[901]), .O(n29458) );
  AO12S U20840 ( .B1(n26080), .B2(n26029), .A1(n26028), .O(n13862) );
  ND2S U20841 ( .I1(n15891), .I2(n26073), .O(n26025) );
  MUX2S U20842 ( .A(n15904), .B(n26073), .S(gray_img[829]), .O(n26026) );
  AO12S U20843 ( .B1(n25936), .B2(n25881), .A1(n25880), .O(n13868) );
  MUX2S U20844 ( .A(n25928), .B(n25929), .S(gray_img[821]), .O(n25878) );
  OA12S U20845 ( .B1(n29831), .B2(n25607), .A1(n25555), .O(n25556) );
  AO12S U20846 ( .B1(n25750), .B2(n25699), .A1(n25698), .O(n13880) );
  ND2S U20847 ( .I1(n15891), .I2(n25744), .O(n25695) );
  MUX2S U20848 ( .A(n25928), .B(n25744), .S(gray_img[805]), .O(n25696) );
  AO12S U20849 ( .B1(n29273), .B2(n29242), .A1(n29241), .O(n13886) );
  MUX2S U20850 ( .A(n30056), .B(n29266), .S(gray_img[797]), .O(n29239) );
  AO12S U20851 ( .B1(n29192), .B2(n29141), .A1(n29140), .O(n13892) );
  ND2S U20852 ( .I1(n27751), .I2(n29186), .O(n29137) );
  AO12S U20853 ( .B1(n29487), .B2(n29436), .A1(n29435), .O(n13904) );
  MUX2S U20854 ( .A(n30044), .B(n29481), .S(gray_img[773]), .O(n29433) );
  ND2S U20855 ( .I1(n28136), .I2(n27934), .O(n27937) );
  OA12S U20856 ( .B1(n29831), .B2(n28139), .A1(n27935), .O(n27936) );
  MUX2S U20857 ( .A(n30005), .B(n28137), .S(gray_img[701]), .O(n27935) );
  AO12S U20858 ( .B1(n28214), .B2(n28105), .A1(n28104), .O(n13932) );
  MUX2S U20859 ( .A(n30005), .B(n28208), .S(gray_img[693]), .O(n28102) );
  AO12S U20860 ( .B1(n28607), .B2(n28436), .A1(n28435), .O(n13939) );
  AO12S U20861 ( .B1(n28588), .B2(n28542), .A1(n28541), .O(n13946) );
  MUX2S U20862 ( .A(n30056), .B(n28581), .S(gray_img[677]), .O(n28539) );
  AO12S U20863 ( .B1(n29350), .B2(n28899), .A1(n28898), .O(n13954) );
  MUX2S U20864 ( .A(n29587), .B(n29344), .S(gray_img[669]), .O(n28896) );
  AO12S U20865 ( .B1(n29040), .B2(n28993), .A1(n28992), .O(n13962) );
  MUX2S U20866 ( .A(n29566), .B(n29033), .S(gray_img[661]), .O(n28990) );
  ND2S U20867 ( .I1(n26445), .I2(n29033), .O(n28989) );
  AO12S U20868 ( .B1(n29904), .B2(n29863), .A1(n29862), .O(n13971) );
  ND2S U20869 ( .I1(n27751), .I2(n29898), .O(n29859) );
  MUX2S U20870 ( .A(n29587), .B(n29898), .S(gray_img[653]), .O(n29860) );
  ND2S U20871 ( .I1(n29993), .I2(n29686), .O(n29689) );
  OA12S U20872 ( .B1(n29831), .B2(n29996), .A1(n29687), .O(n29688) );
  MUX2S U20873 ( .A(n15904), .B(n29994), .S(gray_img[645]), .O(n29687) );
  ND2S U20874 ( .I1(n23492), .I2(n23340), .O(n23343) );
  MUX2S U20875 ( .A(n30050), .B(n23493), .S(gray_img[573]), .O(n23341) );
  AO12S U20876 ( .B1(n28128), .B2(n28074), .A1(n28073), .O(n14014) );
  MUX2S U20877 ( .A(n30050), .B(n28121), .S(gray_img[565]), .O(n28071) );
  AO12S U20878 ( .B1(n28459), .B2(n28405), .A1(n28404), .O(n14023) );
  MUX2S U20879 ( .A(n29032), .B(n28452), .S(gray_img[557]), .O(n28402) );
  ND2S U20880 ( .I1(n28671), .I2(n28561), .O(n28564) );
  OA12S U20881 ( .B1(n29831), .B2(n28674), .A1(n28562), .O(n28563) );
  MUX2S U20882 ( .A(n15904), .B(n28672), .S(gray_img[549]), .O(n28562) );
  AO12S U20883 ( .B1(n28950), .B2(n28904), .A1(n28903), .O(n14041) );
  MUX2S U20884 ( .A(n30056), .B(n28943), .S(gray_img[541]), .O(n28901) );
  ND2S U20885 ( .I1(n29043), .I2(n29017), .O(n29020) );
  MUX2S U20886 ( .A(n30050), .B(n29044), .S(gray_img[533]), .O(n29018) );
  OA12S U20887 ( .B1(n29831), .B2(n29883), .A1(n29830), .O(n29832) );
  MUX2S U20888 ( .A(n30005), .B(n29881), .S(gray_img[525]), .O(n29830) );
  OA12S U20889 ( .B1(n29831), .B2(n29742), .A1(n29712), .O(n29713) );
  MUX2S U20890 ( .A(n15904), .B(n29740), .S(gray_img[517]), .O(n29712) );
  AO12S U20891 ( .B1(n26473), .B2(n26421), .A1(n26420), .O(n14093) );
  ND2S U20892 ( .I1(n26445), .I2(n26466), .O(n26417) );
  MUX2S U20893 ( .A(n15904), .B(n26466), .S(gray_img[445]), .O(n26418) );
  AO12S U20894 ( .B1(n27840), .B2(n26276), .A1(n26275), .O(n14102) );
  ND2S U20895 ( .I1(n15891), .I2(n27834), .O(n26272) );
  MUX2S U20896 ( .A(n15904), .B(n27834), .S(gray_img[437]), .O(n26273) );
  ND2S U20897 ( .I1(n23121), .I2(n23110), .O(n23113) );
  MUX2S U20898 ( .A(n29566), .B(n25151), .S(gray_img[429]), .O(n23111) );
  OA12S U20899 ( .B1(n29831), .B2(n27224), .A1(n23003), .O(n23007) );
  ND2S U20900 ( .I1(n27226), .I2(n23005), .O(n23006) );
  MUX2S U20901 ( .A(n30056), .B(n27222), .S(gray_img[421]), .O(n23003) );
  AO12S U20902 ( .B1(n26489), .B2(n26450), .A1(n26449), .O(n14137) );
  MUX2S U20903 ( .A(n15904), .B(n26483), .S(gray_img[317]), .O(n26447) );
  ND2S U20904 ( .I1(n26327), .I2(n26298), .O(n26299) );
  OA12S U20905 ( .B1(n29831), .B2(n26324), .A1(n26297), .O(n26300) );
  MUX2S U20906 ( .A(n15904), .B(n26322), .S(gray_img[309]), .O(n26297) );
  AO12S U20907 ( .B1(n27121), .B2(n27087), .A1(n27086), .O(n14155) );
  MUX2S U20908 ( .A(n29566), .B(n27114), .S(gray_img[301]), .O(n27084) );
  ND2S U20909 ( .I1(n27751), .I2(n27114), .O(n27083) );
  OA12S U20910 ( .B1(n29831), .B2(n27254), .A1(n27203), .O(n27204) );
  ND2S U20911 ( .I1(n27251), .I2(n27202), .O(n27205) );
  MUX2S U20912 ( .A(n15904), .B(n27252), .S(gray_img[293]), .O(n27203) );
  AO12S U20913 ( .B1(n27692), .B2(n27641), .A1(n27640), .O(n14181) );
  ND2S U20914 ( .I1(n27751), .I2(n27685), .O(n27637) );
  MUX2S U20915 ( .A(n30050), .B(n27685), .S(gray_img[189]), .O(n27638) );
  AO12S U20916 ( .B1(n27785), .B2(n27496), .A1(n27495), .O(n14190) );
  ND2S U20917 ( .I1(n15891), .I2(n27779), .O(n27492) );
  MUX2S U20918 ( .A(n15904), .B(n27779), .S(gray_img[181]), .O(n27493) );
  AO12S U20919 ( .B1(n26939), .B2(n26908), .A1(n26907), .O(n14208) );
  MUX2S U20920 ( .A(n29032), .B(n26932), .S(gray_img[165]), .O(n26905) );
  ND2S U20921 ( .I1(n26828), .I2(n26932), .O(n26904) );
  AO12S U20922 ( .B1(n27708), .B2(n27669), .A1(n27668), .O(n14225) );
  MUX2S U20923 ( .A(n15904), .B(n27702), .S(gray_img[61]), .O(n27666) );
  AO12S U20924 ( .B1(n27556), .B2(n27522), .A1(n27521), .O(n14234) );
  MUX2S U20925 ( .A(n29032), .B(n27550), .S(gray_img[53]), .O(n27519) );
  ND2S U20926 ( .I1(n26445), .I2(n27550), .O(n27518) );
  AO12S U20927 ( .B1(n26849), .B2(n26833), .A1(n26832), .O(n14243) );
  MUX2S U20928 ( .A(n29032), .B(n26842), .S(gray_img[45]), .O(n26830) );
  AO12S U20929 ( .B1(n26931), .B2(n26888), .A1(n26887), .O(n14252) );
  ND2S U20930 ( .I1(n27751), .I2(n26924), .O(n26884) );
  MUX2S U20931 ( .A(n30056), .B(n26924), .S(gray_img[37]), .O(n26885) );
  AO12S U20932 ( .B1(n27751), .B2(n25836), .A1(n25826), .O(n15080) );
  MUX2S U20933 ( .A(n28534), .B(n25834), .S(gray_img[2021]), .O(n25826) );
  AO12S U20934 ( .B1(n26445), .B2(n25473), .A1(n25462), .O(n15081) );
  MUX2S U20935 ( .A(n28534), .B(n25471), .S(gray_img[2013]), .O(n25462) );
  AO12S U20936 ( .B1(n27751), .B2(n25761), .A1(n25449), .O(n15082) );
  AO12S U20937 ( .B1(n15891), .B2(n28803), .A1(n25625), .O(n15083) );
  MUX2S U20938 ( .A(n29566), .B(n20746), .S(gray_img[1981]), .O(n18856) );
  MUX2S U20939 ( .A(n29597), .B(n20849), .S(gray_img[1973]), .O(n18692) );
  MUX2S U20940 ( .A(n29587), .B(n19970), .S(gray_img[1949]), .O(n18634) );
  MUX2S U20941 ( .A(n30056), .B(n20389), .S(gray_img[1941]), .O(n18901) );
  MUX2S U20942 ( .A(n30044), .B(n20424), .S(gray_img[1933]), .O(n18810) );
  MUX2S U20943 ( .A(n20842), .B(n20373), .S(gray_img[1925]), .O(n18880) );
  MUX2S U20944 ( .A(n30050), .B(n20430), .S(gray_img[1917]), .O(n18750) );
  MUX2S U20945 ( .A(n29587), .B(n20063), .S(gray_img[1909]), .O(n18530) );
  MUX2S U20946 ( .A(n30056), .B(n20544), .S(gray_img[1901]), .O(n18952) );
  AO12S U20947 ( .B1(n15891), .B2(n25832), .A1(n25821), .O(n15096) );
  MUX2S U20948 ( .A(n27447), .B(n25830), .S(gray_img[1893]), .O(n25821) );
  AO12S U20949 ( .B1(n15891), .B2(n25477), .A1(n25467), .O(n15097) );
  MUX2S U20950 ( .A(n27447), .B(n25475), .S(gray_img[1885]), .O(n25467) );
  AO12S U20951 ( .B1(n15891), .B2(n25460), .A1(n25450), .O(n15098) );
  MUX2S U20952 ( .A(n27447), .B(n25458), .S(gray_img[1877]), .O(n25450) );
  AO12S U20953 ( .B1(n26828), .B2(n25631), .A1(n25620), .O(n15099) );
  MUX2S U20954 ( .A(n29597), .B(n20504), .S(gray_img[1861]), .O(n18983) );
  MUX2S U20955 ( .A(n29566), .B(n20740), .S(gray_img[1853]), .O(n18852) );
  MUX2S U20956 ( .A(n29597), .B(n20862), .S(gray_img[1845]), .O(n18682) );
  MUX2S U20957 ( .A(n29587), .B(n20296), .S(gray_img[1821]), .O(n18628) );
  MUX2S U20958 ( .A(n29566), .B(n20354), .S(gray_img[1813]), .O(n20337) );
  MUX2S U20959 ( .A(n30050), .B(n20319), .S(gray_img[1805]), .O(n18814) );
  MUX2S U20960 ( .A(n20842), .B(n20547), .S(gray_img[1789]), .O(n18805) );
  MUX2S U20961 ( .A(n30044), .B(n20449), .S(gray_img[1773]), .O(n18955) );
  AO12S U20962 ( .B1(n15891), .B2(n25778), .A1(n25767), .O(n15112) );
  MUX2S U20963 ( .A(n15889), .B(n25776), .S(gray_img[1765]), .O(n25767) );
  AO12S U20964 ( .B1(n26445), .B2(n25510), .A1(n25499), .O(n15113) );
  MUX2S U20965 ( .A(n27447), .B(n25508), .S(gray_img[1757]), .O(n25499) );
  AO12S U20966 ( .B1(n26828), .B2(n25498), .A1(n25488), .O(n15114) );
  MUX2S U20967 ( .A(n28534), .B(n25496), .S(gray_img[1749]), .O(n25488) );
  AO12S U20968 ( .B1(n15891), .B2(n25649), .A1(n25638), .O(n15115) );
  MUX2S U20969 ( .A(n29597), .B(n19955), .S(gray_img[1733]), .O(n18986) );
  MUX2S U20970 ( .A(n30044), .B(n20737), .S(gray_img[1725]), .O(n18834) );
  MUX2S U20971 ( .A(n30056), .B(n20846), .S(gray_img[1717]), .O(n18685) );
  MUX2S U20972 ( .A(n30050), .B(n20827), .S(gray_img[1709]), .O(n18759) );
  MUX2S U20973 ( .A(n30056), .B(n20787), .S(gray_img[1701]), .O(n18520) );
  MUX2S U20974 ( .A(n29566), .B(n20605), .S(gray_img[1685]), .O(n18895) );
  MUX2S U20975 ( .A(n29566), .B(n20531), .S(gray_img[1677]), .O(n18714) );
  MUX2S U20976 ( .A(n29566), .B(n20583), .S(gray_img[1669]), .O(n18847) );
  MUX2S U20977 ( .A(n29587), .B(n20509), .S(gray_img[1661]), .O(n18764) );
  MUX2S U20978 ( .A(n29566), .B(n20525), .S(gray_img[1653]), .O(n18547) );
  AO12S U20979 ( .B1(n15891), .B2(n25899), .A1(n25772), .O(n15128) );
  AO12S U20980 ( .B1(n15891), .B2(n25576), .A1(n25504), .O(n15129) );
  AO12S U20981 ( .B1(n27751), .B2(n25494), .A1(n25483), .O(n15130) );
  AO12S U20982 ( .B1(n15891), .B2(n25653), .A1(n25643), .O(n15131) );
  MUX2S U20983 ( .A(n28534), .B(n25651), .S(gray_img[1613]), .O(n25643) );
  MUX2S U20984 ( .A(n15904), .B(n20528), .S(gray_img[1605]), .O(n18981) );
  MUX2S U20985 ( .A(n30056), .B(n20731), .S(gray_img[1597]), .O(n18837) );
  MUX2S U20986 ( .A(n20830), .B(n20839), .S(gray_img[1589]), .O(n18665) );
  MUX2S U20987 ( .A(n30050), .B(n20395), .S(gray_img[1581]), .O(n18762) );
  MUX2S U20988 ( .A(n30056), .B(n20824), .S(gray_img[1573]), .O(n18523) );
  MUX2S U20989 ( .A(n29587), .B(n20602), .S(gray_img[1557]), .O(n18898) );
  MUX2S U20990 ( .A(n29587), .B(n20550), .S(gray_img[1549]), .O(n18709) );
  MUX2S U20991 ( .A(n29597), .B(n20881), .S(gray_img[1541]), .O(n20872) );
  MUX2S U20992 ( .A(n30050), .B(n20556), .S(gray_img[1533]), .O(n18745) );
  MUX2S U20993 ( .A(n20808), .B(n20512), .S(gray_img[1525]), .O(n18817) );
  MUX2S U20994 ( .A(n30056), .B(n20440), .S(gray_img[1517]), .O(n18975) );
  AO12S U20995 ( .B1(n26445), .B2(n27971), .A1(n27961), .O(n15144) );
  MUX2S U20996 ( .A(n28534), .B(n27969), .S(gray_img[1509]), .O(n27961) );
  AO12S U20997 ( .B1(n26828), .B2(n28355), .A1(n28344), .O(n15145) );
  MUX2S U20998 ( .A(n28534), .B(n28353), .S(gray_img[1501]), .O(n28344) );
  AO12S U20999 ( .B1(n15891), .B2(n28342), .A1(n28331), .O(n15146) );
  MUX2S U21000 ( .A(n27447), .B(n28340), .S(gray_img[1493]), .O(n28331) );
  AO12S U21001 ( .B1(n15891), .B2(n28560), .A1(n28528), .O(n15147) );
  MUX2S U21002 ( .A(n15889), .B(n28558), .S(gray_img[1485]), .O(n28528) );
  MUX2S U21003 ( .A(n15904), .B(n20684), .S(gray_img[1477]), .O(n18999) );
  MUX2S U21004 ( .A(n20830), .B(n20709), .S(gray_img[1469]), .O(n18827) );
  MUX2S U21005 ( .A(n30056), .B(n20821), .S(gray_img[1461]), .O(n18668) );
  MUX2S U21006 ( .A(n30044), .B(n20811), .S(gray_img[1445]), .O(n18575) );
  MUX2S U21007 ( .A(n30044), .B(n20293), .S(gray_img[1437]), .O(n18601) );
  MUX2S U21008 ( .A(n20842), .B(n20193), .S(gray_img[1429]), .O(n18887) );
  MUX2S U21009 ( .A(n20842), .B(n20035), .S(gray_img[1421]), .O(n18703) );
  MUX2S U21010 ( .A(n30044), .B(n20571), .S(gray_img[1405]), .O(n18748) );
  MUX2S U21011 ( .A(n20808), .B(n20517), .S(gray_img[1397]), .O(n18831) );
  MUX2S U21012 ( .A(n30050), .B(n20722), .S(gray_img[1389]), .O(n18969) );
  ND2S U21013 ( .I1(n27447), .I2(n27993), .O(n27959) );
  AO12S U21014 ( .B1(n15891), .B2(n28359), .A1(n28349), .O(n15161) );
  MUX2S U21015 ( .A(n27447), .B(n28357), .S(gray_img[1373]), .O(n28349) );
  AO12S U21016 ( .B1(n27751), .B2(n28596), .A1(n28336), .O(n15162) );
  MUX2S U21017 ( .A(n28534), .B(n28594), .S(gray_img[1365]), .O(n28336) );
  AO12S U21018 ( .B1(n15891), .B2(n28536), .A1(n28523), .O(n15163) );
  MUX2S U21019 ( .A(n28534), .B(n28533), .S(gray_img[1357]), .O(n28523) );
  MUX2S U21020 ( .A(n15904), .B(n20734), .S(gray_img[1349]), .O(n19005) );
  MUX2S U21021 ( .A(n20830), .B(n20695), .S(gray_img[1341]), .O(n18824) );
  MUX2S U21022 ( .A(n30044), .B(n20833), .S(gray_img[1333]), .O(n18676) );
  MUX2S U21023 ( .A(n29566), .B(n20836), .S(gray_img[1325]), .O(n18777) );
  MUX2S U21024 ( .A(n30044), .B(n20362), .S(gray_img[1301]), .O(n18890) );
  MUX2S U21025 ( .A(n20842), .B(n20427), .S(gray_img[1293]), .O(n18706) );
  MUX2S U21026 ( .A(n15904), .B(n20392), .S(gray_img[1285]), .O(n18863) );
  MUX2S U21027 ( .A(n20808), .B(n20655), .S(gray_img[1277]), .O(n18799) );
  MUX2S U21028 ( .A(n20808), .B(n20725), .S(gray_img[1269]), .O(n18592) );
  MUX2S U21029 ( .A(n30044), .B(n20719), .S(gray_img[1261]), .O(n18971) );
  AO12S U21030 ( .B1(n15891), .B2(n28031), .A1(n28024), .O(n15176) );
  MUX2S U21031 ( .A(n28534), .B(n28029), .S(gray_img[1253]), .O(n28024) );
  AO12S U21032 ( .B1(n15891), .B2(n28288), .A1(n28278), .O(n15177) );
  MUX2S U21033 ( .A(n28534), .B(n28286), .S(gray_img[1245]), .O(n28278) );
  AO12S U21034 ( .B1(n15891), .B2(n28271), .A1(n28260), .O(n15178) );
  AO12S U21035 ( .B1(n27751), .B2(n28475), .A1(n28465), .O(n15179) );
  MUX2S U21036 ( .A(n28534), .B(n28473), .S(gray_img[1229]), .O(n28465) );
  MUX2S U21037 ( .A(n29587), .B(n20702), .S(gray_img[1221]), .O(n19003) );
  ND2S U21038 ( .I1(n19741), .I2(n19740), .O(n15181) );
  MUX2S U21039 ( .A(n30044), .B(n20757), .S(gray_img[1213]), .O(n19740) );
  MUX2S U21040 ( .A(n30044), .B(n20857), .S(gray_img[1205]), .O(n18671) );
  MUX2S U21041 ( .A(n29587), .B(n20435), .S(gray_img[1197]), .O(n19670) );
  MUX2S U21042 ( .A(n29566), .B(n20379), .S(gray_img[1189]), .O(n18557) );
  MUX2S U21043 ( .A(n29597), .B(n20159), .S(gray_img[1181]), .O(n18613) );
  MUX2S U21044 ( .A(n30056), .B(n20316), .S(gray_img[1173]), .O(n19760) );
  MUX2S U21045 ( .A(n29587), .B(n20553), .S(gray_img[1165]), .O(n18719) );
  MUX2S U21046 ( .A(n30005), .B(n20240), .S(gray_img[1157]), .O(n19702) );
  MUX2S U21047 ( .A(n30050), .B(n20716), .S(gray_img[1149]), .O(n18803) );
  MUX2S U21048 ( .A(n20808), .B(n20124), .S(gray_img[1141]), .O(n18594) );
  MUX2S U21049 ( .A(n30044), .B(n20728), .S(gray_img[1133]), .O(n18958) );
  AO12S U21050 ( .B1(n15891), .B2(n28092), .A1(n28019), .O(n15192) );
  MUX2S U21051 ( .A(n28534), .B(n28090), .S(gray_img[1125]), .O(n28019) );
  AO12S U21052 ( .B1(n15891), .B2(n28284), .A1(n28273), .O(n15193) );
  AO12S U21053 ( .B1(n15891), .B2(n28423), .A1(n28265), .O(n15194) );
  MUX2S U21054 ( .A(n27447), .B(n28421), .S(gray_img[1109]), .O(n28265) );
  AO12S U21055 ( .B1(n15891), .B2(n28480), .A1(n28467), .O(n15195) );
  MUX2S U21056 ( .A(n27447), .B(n28478), .S(gray_img[1101]), .O(n28467) );
  MUX2S U21057 ( .A(n30050), .B(n20743), .S(gray_img[1093]), .O(n18996) );
  ND2S U21058 ( .I1(n19743), .I2(n19742), .O(n15197) );
  MUX2S U21059 ( .A(n30056), .B(n20760), .S(gray_img[1085]), .O(n19742) );
  MUX2S U21060 ( .A(n30044), .B(n20854), .S(gray_img[1077]), .O(n18679) );
  MUX2S U21061 ( .A(n30044), .B(n20611), .S(gray_img[1069]), .O(n19665) );
  MUX2S U21062 ( .A(n29587), .B(n20368), .S(gray_img[1061]), .O(n18555) );
  MUX2S U21063 ( .A(n30044), .B(n20184), .S(gray_img[1053]), .O(n18618) );
  ND2S U21064 ( .I1(n19777), .I2(n19776), .O(n15202) );
  MUX2S U21065 ( .A(n29597), .B(n20255), .S(gray_img[1045]), .O(n19776) );
  MUX2S U21066 ( .A(n29587), .B(n20235), .S(gray_img[1037]), .O(n19418) );
  MUX2S U21067 ( .A(n15904), .B(n20099), .S(gray_img[1021]), .O(n18661) );
  MUX2S U21068 ( .A(n20808), .B(n20562), .S(gray_img[1013]), .O(n18540) );
  AO12S U21069 ( .B1(n26828), .B2(n27829), .A1(n26218), .O(n15208) );
  AO12S U21070 ( .B1(n15891), .B2(n27081), .A1(n27070), .O(n15209) );
  AO12S U21071 ( .B1(n15891), .B2(n27065), .A1(n27054), .O(n15210) );
  MUX2S U21072 ( .A(n29587), .B(n20580), .S(gray_img[965]), .O(n18931) );
  MUX2S U21073 ( .A(n30044), .B(n20452), .S(gray_img[893]), .O(n18655) );
  MUX2S U21074 ( .A(n15904), .B(n20559), .S(gray_img[885]), .O(n18545) );
  AO12S U21075 ( .B1(n15891), .B2(n26224), .A1(n26213), .O(n15216) );
  AO12S U21076 ( .B1(n15891), .B2(n30065), .A1(n27075), .O(n15217) );
  MUX2S U21077 ( .A(n15889), .B(n30063), .S(gray_img[861]), .O(n27075) );
  AO12S U21078 ( .B1(n26445), .B2(n27069), .A1(n27059), .O(n15218) );
  ND2S U21079 ( .I1(n19923), .I2(n19922), .O(n15220) );
  MUX2S U21080 ( .A(n29587), .B(n20634), .S(gray_img[837]), .O(n19922) );
  MUX2S U21081 ( .A(n25928), .B(n20568), .S(gray_img[765]), .O(n18649) );
  MUX2S U21082 ( .A(n30005), .B(n20054), .S(gray_img[757]), .O(n18550) );
  AO12S U21083 ( .B1(n15891), .B2(n26155), .A1(n26145), .O(n15224) );
  AO12S U21084 ( .B1(n15891), .B2(n26996), .A1(n26985), .O(n15225) );
  MUX2S U21085 ( .A(n27447), .B(n26994), .S(gray_img[733]), .O(n26985) );
  AO12S U21086 ( .B1(n15891), .B2(n27009), .A1(n26998), .O(n15226) );
  AO12S U21087 ( .B1(n15891), .B2(n27243), .A1(n27127), .O(n15227) );
  MUX2S U21088 ( .A(n28534), .B(n27241), .S(gray_img[717]), .O(n27127) );
  ND2S U21089 ( .I1(n19867), .I2(n19866), .O(n15228) );
  MUX2S U21090 ( .A(n15904), .B(n20623), .S(gray_img[709]), .O(n19866) );
  MUX2S U21091 ( .A(n29597), .B(n20565), .S(gray_img[637]), .O(n18658) );
  MUX2S U21092 ( .A(n30050), .B(n20534), .S(gray_img[629]), .O(n18535) );
  ND2S U21093 ( .I1(n19839), .I2(n19838), .O(n15231) );
  AO12S U21094 ( .B1(n15891), .B2(n26160), .A1(n26157), .O(n15232) );
  AO12S U21095 ( .B1(n15891), .B2(n27105), .A1(n26990), .O(n15233) );
  AO12S U21096 ( .B1(n15891), .B2(n27013), .A1(n27003), .O(n15234) );
  AO12S U21097 ( .B1(n15891), .B2(n27133), .A1(n27122), .O(n15235) );
  MUX2S U21098 ( .A(n15889), .B(n27131), .S(gray_img[589]), .O(n27122) );
  MUX2S U21099 ( .A(n29597), .B(n20591), .S(gray_img[581]), .O(n18925) );
  MUX2S U21100 ( .A(n20830), .B(n20472), .S(gray_img[509]), .O(n18807) );
  MUX2S U21101 ( .A(n30056), .B(n20477), .S(gray_img[501]), .O(n18528) );
  MUX2S U21102 ( .A(n29597), .B(n20480), .S(gray_img[493]), .O(n19812) );
  AO12S U21103 ( .B1(n15891), .B2(n27774), .A1(n27442), .O(n15240) );
  AO12S U21104 ( .B1(n15891), .B2(n27352), .A1(n26753), .O(n15241) );
  MUX2S U21105 ( .A(n28534), .B(n27350), .S(gray_img[477]), .O(n26753) );
  AO12S U21106 ( .B1(n15891), .B2(n26747), .A1(n26736), .O(n15242) );
  MUX2S U21107 ( .A(n27447), .B(n26745), .S(gray_img[469]), .O(n26736) );
  AO12S U21108 ( .B1(n15891), .B2(n26942), .A1(n26855), .O(n15243) );
  MUX2S U21109 ( .A(n27447), .B(n26940), .S(gray_img[461]), .O(n26855) );
  ND2S U21110 ( .I1(n19876), .I2(n19875), .O(n15244) );
  MUX2S U21111 ( .A(n15904), .B(n20486), .S(gray_img[381]), .O(n18652) );
  MUX2S U21112 ( .A(n30044), .B(n20522), .S(gray_img[373]), .O(n18524) );
  MUX2S U21113 ( .A(n30050), .B(n20491), .S(gray_img[365]), .O(n19801) );
  AO12S U21114 ( .B1(n15891), .B2(n27449), .A1(n27437), .O(n15248) );
  MUX2S U21115 ( .A(n15889), .B(n27446), .S(gray_img[357]), .O(n27437) );
  AO12S U21116 ( .B1(n15891), .B2(n26759), .A1(n26748), .O(n15249) );
  AO12S U21117 ( .B1(n15891), .B2(n26743), .A1(n26732), .O(n15250) );
  MUX2S U21118 ( .A(n27447), .B(n26741), .S(gray_img[341]), .O(n26732) );
  AO12S U21119 ( .B1(n15891), .B2(n26861), .A1(n26850), .O(n15251) );
  MUX2S U21120 ( .A(n29597), .B(n20496), .S(gray_img[253]), .O(n18687) );
  ND2S U21121 ( .I1(n19737), .I2(n19736), .O(n15254) );
  MUX2S U21122 ( .A(n30044), .B(n20260), .S(gray_img[245]), .O(n19736) );
  AO12S U21123 ( .B1(n15891), .B2(n27390), .A1(n27379), .O(n15256) );
  MUX2S U21124 ( .A(n15889), .B(n27388), .S(gray_img[229]), .O(n27379) );
  AO12S U21125 ( .B1(n15891), .B2(n26726), .A1(n26703), .O(n15257) );
  AO12S U21126 ( .B1(n15891), .B2(n26841), .A1(n26716), .O(n15258) );
  AO12S U21127 ( .B1(n26445), .B2(n26883), .A1(n26873), .O(n15259) );
  ND2S U21128 ( .I1(n19899), .I2(n19898), .O(n15260) );
  MUX2S U21129 ( .A(n15904), .B(n20631), .S(gray_img[197]), .O(n19898) );
  MUX2S U21130 ( .A(n29566), .B(n20082), .S(gray_img[125]), .O(n18644) );
  ND2S U21131 ( .I1(n19725), .I2(n19724), .O(n15262) );
  MUX2S U21132 ( .A(n30044), .B(n20499), .S(gray_img[117]), .O(n19724) );
  MUX2S U21133 ( .A(n20617), .B(n20830), .S(n27402), .O(n19847) );
  AO12S U21134 ( .B1(n15891), .B2(n27545), .A1(n27384), .O(n15264) );
  MUX2S U21135 ( .A(n27447), .B(n27543), .S(gray_img[101]), .O(n27384) );
  AO12S U21136 ( .B1(n15891), .B2(n26709), .A1(n26698), .O(n15265) );
  MUX2S U21137 ( .A(n27447), .B(n26707), .S(gray_img[93]), .O(n26698) );
  MUX2S U21138 ( .A(n15889), .B(n26720), .S(gray_img[85]), .O(n26711) );
  AO12S U21139 ( .B1(n15891), .B2(n26879), .A1(n26868), .O(n15267) );
  MUX2S U21140 ( .A(n27447), .B(n26877), .S(gray_img[77]), .O(n26868) );
  ND2S U21141 ( .I1(n19910), .I2(n19909), .O(n15268) );
  MUX2S U21142 ( .A(n15904), .B(n20628), .S(gray_img[69]), .O(n19909) );
  ND2S U21143 ( .I1(n22961), .I2(n22960), .O(n15810) );
  ND2S U21144 ( .I1(n30120), .I2(n23468), .O(n23471) );
  AO12S U21145 ( .B1(n28847), .B2(n28780), .A1(n28779), .O(n15272) );
  ND2S U21146 ( .I1(n28727), .I2(n26135), .O(n26138) );
  AO12S U21147 ( .B1(n28724), .B2(n25983), .A1(n25982), .O(n13614) );
  MUX2S U21148 ( .A(n15904), .B(n28718), .S(gray_img[958]), .O(n25980) );
  AO12S U21149 ( .B1(n26096), .B2(n25876), .A1(n25875), .O(n13615) );
  ND2S U21150 ( .I1(n15890), .I2(n26090), .O(n25872) );
  MUX2S U21151 ( .A(n15904), .B(n26090), .S(gray_img[950]), .O(n25873) );
  ND2S U21152 ( .I1(n28806), .I2(n25762), .O(n25765) );
  MUX2S U21153 ( .A(n29566), .B(n28807), .S(gray_img[406]), .O(n25763) );
  ND2S U21154 ( .I1(n30128), .I2(n18135), .O(n18143) );
  AO12S U21155 ( .B1(n30109), .B2(n29644), .A1(n29643), .O(n13632) );
  MUX2S U21156 ( .A(n15904), .B(n30103), .S(gray_img[390]), .O(n29641) );
  ND2S U21157 ( .I1(n28247), .I2(n28181), .O(n28184) );
  OA12S U21158 ( .B1(n29825), .B2(n28250), .A1(n28182), .O(n28183) );
  MUX2S U21159 ( .A(n30005), .B(n28248), .S(gray_img[286]), .O(n28182) );
  ND2S U21160 ( .I1(n28706), .I2(n28644), .O(n28647) );
  AO12S U21161 ( .B1(n29381), .B2(n29096), .A1(n29095), .O(n13701) );
  MUX2S U21162 ( .A(n30056), .B(n29374), .S(gray_img[270]), .O(n29093) );
  AO12S U21163 ( .B1(n30012), .B2(n29945), .A1(n29944), .O(n13730) );
  MUX2S U21164 ( .A(n30005), .B(n30006), .S(gray_img[262]), .O(n29942) );
  ND2S U21165 ( .I1(n30087), .I2(n27888), .O(n27891) );
  AO12S U21166 ( .B1(n27851), .B2(n26528), .A1(n26527), .O(n13756) );
  MUX2S U21167 ( .A(n29597), .B(n27845), .S(gray_img[158]), .O(n26525) );
  AO12S U21168 ( .B1(n30076), .B2(n27303), .A1(n27302), .O(n13766) );
  MUX2S U21169 ( .A(n15904), .B(n30070), .S(gray_img[150]), .O(n27300) );
  AO12S U21170 ( .B1(n27821), .B2(n27750), .A1(n27749), .O(n13786) );
  MUX2S U21171 ( .A(n30005), .B(n27814), .S(gray_img[30]), .O(n27747) );
  AO12S U21172 ( .B1(n27378), .B2(n26984), .A1(n26983), .O(n13796) );
  MUX2S U21173 ( .A(n30005), .B(n27371), .S(gray_img[22]), .O(n26981) );
  AO12S U21174 ( .B1(n25758), .B2(n25637), .A1(n25636), .O(n13821) );
  ND2S U21175 ( .I1(n15890), .I2(n25751), .O(n25633) );
  MUX2S U21176 ( .A(n30056), .B(n25751), .S(gray_img[934]), .O(n25634) );
  AO12S U21177 ( .B1(n30038), .B2(n29314), .A1(n29313), .O(n15071) );
  MUX2S U21178 ( .A(n30056), .B(n30032), .S(gray_img[398]), .O(n29311) );
  ND2S U21179 ( .I1(n30020), .I2(n26693), .O(n26696) );
  AO12S U21180 ( .B1(n29604), .B2(n29530), .A1(n29529), .O(n13834) );
  MUX2S U21181 ( .A(n30044), .B(n29598), .S(gray_img[910]), .O(n29527) );
  ND2S U21182 ( .I1(n30098), .I2(n29426), .O(n29430) );
  AO12S U21183 ( .B1(n26080), .B2(n26024), .A1(n26023), .O(n13861) );
  MUX2S U21184 ( .A(n15904), .B(n26073), .S(gray_img[830]), .O(n26021) );
  AO12S U21185 ( .B1(n25936), .B2(n25820), .A1(n25819), .O(n13867) );
  MUX2S U21186 ( .A(n25928), .B(n25929), .S(gray_img[822]), .O(n25817) );
  AO12S U21187 ( .B1(n25750), .B2(n25694), .A1(n25693), .O(n13879) );
  MUX2S U21188 ( .A(n25928), .B(n25744), .S(gray_img[806]), .O(n25691) );
  ND2S U21189 ( .I1(n29273), .I2(n29233), .O(n29236) );
  AO12S U21190 ( .B1(n29192), .B2(n29136), .A1(n29135), .O(n13891) );
  ND2S U21191 ( .I1(n29579), .I2(n26570), .O(n26573) );
  AO12S U21192 ( .B1(n29487), .B2(n26616), .A1(n26615), .O(n13903) );
  MUX2S U21193 ( .A(n30056), .B(n29481), .S(gray_img[774]), .O(n26613) );
  ND2S U21194 ( .I1(n28136), .I2(n27929), .O(n27932) );
  OA12S U21195 ( .B1(n29825), .B2(n28139), .A1(n27930), .O(n27931) );
  MUX2S U21196 ( .A(n30005), .B(n28137), .S(gray_img[702]), .O(n27930) );
  AO12S U21197 ( .B1(n28214), .B2(n28018), .A1(n28017), .O(n13931) );
  MUX2S U21198 ( .A(n30005), .B(n28208), .S(gray_img[694]), .O(n28015) );
  AO12S U21199 ( .B1(n28607), .B2(n28400), .A1(n28399), .O(n13938) );
  ND2S U21200 ( .I1(n29350), .I2(n18093), .O(n18100) );
  AO12S U21201 ( .B1(n29040), .B2(n28988), .A1(n28987), .O(n13961) );
  MUX2S U21202 ( .A(n29587), .B(n29033), .S(gray_img[662]), .O(n28985) );
  AO12S U21203 ( .B1(n29904), .B2(n29788), .A1(n29787), .O(n13970) );
  MUX2S U21204 ( .A(n29566), .B(n29898), .S(gray_img[654]), .O(n29785) );
  ND2S U21205 ( .I1(n29993), .I2(n29681), .O(n29684) );
  OA12S U21206 ( .B1(n29825), .B2(n29996), .A1(n29682), .O(n29683) );
  MUX2S U21207 ( .A(n15904), .B(n29994), .S(gray_img[646]), .O(n29682) );
  ND2S U21208 ( .I1(n23492), .I2(n23350), .O(n23353) );
  MUX2S U21209 ( .A(n30044), .B(n23493), .S(gray_img[574]), .O(n23351) );
  AO12S U21210 ( .B1(n28128), .B2(n28069), .A1(n28068), .O(n14013) );
  MUX2S U21211 ( .A(n30005), .B(n28121), .S(gray_img[566]), .O(n28066) );
  AO12S U21212 ( .B1(n28459), .B2(n28330), .A1(n28329), .O(n14022) );
  MUX2S U21213 ( .A(n29032), .B(n28452), .S(gray_img[558]), .O(n28327) );
  ND2S U21214 ( .I1(n28671), .I2(n28518), .O(n28521) );
  OA12S U21215 ( .B1(n29825), .B2(n28674), .A1(n28519), .O(n28520) );
  MUX2S U21216 ( .A(n15904), .B(n28672), .S(gray_img[550]), .O(n28519) );
  AO12S U21217 ( .B1(n28950), .B2(n28894), .A1(n28893), .O(n14040) );
  MUX2S U21218 ( .A(n30050), .B(n28943), .S(gray_img[542]), .O(n28891) );
  ND2S U21219 ( .I1(n29043), .I2(n26140), .O(n26143) );
  MUX2S U21220 ( .A(n30050), .B(n29044), .S(gray_img[534]), .O(n26141) );
  OA12S U21221 ( .B1(n29825), .B2(n29883), .A1(n29824), .O(n29826) );
  MUX2S U21222 ( .A(n30005), .B(n29881), .S(gray_img[526]), .O(n29824) );
  ND2S U21223 ( .I1(n29739), .I2(n26651), .O(n26654) );
  AO12S U21224 ( .B1(n26473), .B2(n26416), .A1(n26415), .O(n14092) );
  MUX2S U21225 ( .A(n29566), .B(n26466), .S(gray_img[446]), .O(n26413) );
  AO12S U21226 ( .B1(n27840), .B2(n26271), .A1(n26270), .O(n14101) );
  MUX2S U21227 ( .A(n30050), .B(n27834), .S(gray_img[438]), .O(n26268) );
  ND2S U21228 ( .I1(n23121), .I2(n23115), .O(n23118) );
  OA12S U21229 ( .B1(n29825), .B2(n27224), .A1(n27192), .O(n27195) );
  ND2S U21230 ( .I1(n27226), .I2(n27193), .O(n27194) );
  MUX2S U21231 ( .A(n30056), .B(n27222), .S(gray_img[422]), .O(n27192) );
  ND2S U21232 ( .I1(n26489), .I2(n26370), .O(n26373) );
  ND2S U21233 ( .I1(n26327), .I2(n26209), .O(n26210) );
  OA12S U21234 ( .B1(n29825), .B2(n26324), .A1(n26206), .O(n26211) );
  AO12S U21235 ( .B1(n27121), .B2(n27053), .A1(n27052), .O(n14154) );
  MUX2S U21236 ( .A(n29597), .B(n27114), .S(gray_img[302]), .O(n27050) );
  OA12S U21237 ( .B1(n29825), .B2(n27254), .A1(n27171), .O(n27172) );
  ND2S U21238 ( .I1(n27251), .I2(n27170), .O(n27173) );
  MUX2S U21239 ( .A(n15904), .B(n27252), .S(gray_img[294]), .O(n27171) );
  AO12S U21240 ( .B1(n27692), .B2(n27636), .A1(n27635), .O(n14180) );
  MUX2S U21241 ( .A(n30044), .B(n27685), .S(gray_img[190]), .O(n27633) );
  AO12S U21242 ( .B1(n27785), .B2(n27491), .A1(n27490), .O(n14189) );
  MUX2S U21243 ( .A(n15904), .B(n27779), .S(gray_img[182]), .O(n27488) );
  OA12S U21244 ( .B1(n29825), .B2(n27358), .A1(n26799), .O(n26800) );
  MUX2S U21245 ( .A(n29587), .B(n27356), .S(gray_img[174]), .O(n26799) );
  AO12S U21246 ( .B1(n26939), .B2(n26867), .A1(n26866), .O(n14207) );
  MUX2S U21247 ( .A(n29032), .B(n26932), .S(gray_img[166]), .O(n26864) );
  AO12S U21248 ( .B1(n27708), .B2(n27598), .A1(n27597), .O(n14224) );
  MUX2S U21249 ( .A(n15904), .B(n27702), .S(gray_img[62]), .O(n27595) );
  AO12S U21250 ( .B1(n27556), .B2(n27436), .A1(n27435), .O(n14233) );
  MUX2S U21251 ( .A(n29032), .B(n27550), .S(gray_img[54]), .O(n27433) );
  AO12S U21252 ( .B1(n26849), .B2(n26731), .A1(n26730), .O(n14242) );
  MUX2S U21253 ( .A(n29032), .B(n26842), .S(gray_img[46]), .O(n26728) );
  ND2S U21254 ( .I1(n26931), .I2(n23632), .O(n23635) );
  AO12S U21255 ( .B1(n25619), .B2(n25482), .A1(n25481), .O(n15270) );
  MUX2S U21256 ( .A(n30050), .B(n25612), .S(gray_img[942]), .O(n25479) );
  ND2S U21257 ( .I1(n20417), .I2(n20416), .O(n15275) );
  MUX2S U21258 ( .A(n30005), .B(n20608), .S(gray_img[2030]), .O(n20416) );
  AO12S U21259 ( .B1(n25444), .B2(n25836), .A1(n25439), .O(n15276) );
  MUX2S U21260 ( .A(n28534), .B(n25834), .S(gray_img[2022]), .O(n25439) );
  AO12S U21261 ( .B1(n25448), .B2(n25473), .A1(n25381), .O(n15277) );
  ND2S U21262 ( .I1(n15889), .I2(n25403), .O(n25404) );
  AO12S U21263 ( .B1(n25444), .B2(n28803), .A1(n25414), .O(n15279) );
  MUX2S U21264 ( .A(n27447), .B(n28801), .S(gray_img[1998]), .O(n25414) );
  ND2S U21265 ( .I1(n18940), .I2(n18939), .O(n15280) );
  MUX2S U21266 ( .A(n29597), .B(n20209), .S(gray_img[1990]), .O(n18940) );
  ND2S U21267 ( .I1(n20419), .I2(n20418), .O(n15281) );
  MUX2S U21268 ( .A(n29566), .B(n20746), .S(gray_img[1982]), .O(n20418) );
  ND2S U21269 ( .I1(n20358), .I2(n20357), .O(n15282) );
  MUX2S U21270 ( .A(n29597), .B(n20849), .S(gray_img[1974]), .O(n20358) );
  ND2S U21271 ( .I1(n20006), .I2(n20005), .O(n15283) );
  ND2S U21272 ( .I1(n20347), .I2(n20346), .O(n15284) );
  MUX2S U21273 ( .A(n30056), .B(n19970), .S(gray_img[1950]), .O(n18610) );
  ND2S U21274 ( .I1(n20391), .I2(n20390), .O(n15286) );
  MUX2S U21275 ( .A(n30050), .B(n20389), .S(gray_img[1942]), .O(n20391) );
  ND2S U21276 ( .I1(n20426), .I2(n20425), .O(n15287) );
  MUX2S U21277 ( .A(n30056), .B(n20424), .S(gray_img[1934]), .O(n20425) );
  ND2S U21278 ( .I1(n20375), .I2(n20374), .O(n15288) );
  MUX2S U21279 ( .A(n20842), .B(n20373), .S(gray_img[1926]), .O(n20375) );
  ND2S U21280 ( .I1(n20432), .I2(n20431), .O(n15289) );
  MUX2S U21281 ( .A(n15904), .B(n20430), .S(gray_img[1918]), .O(n20431) );
  ND2S U21282 ( .I1(n20403), .I2(n20402), .O(n15291) );
  MUX2S U21283 ( .A(n30056), .B(n20544), .S(gray_img[1902]), .O(n20402) );
  AO12S U21284 ( .B1(n25448), .B2(n25832), .A1(n25430), .O(n15292) );
  MUX2S U21285 ( .A(n28534), .B(n25830), .S(gray_img[1894]), .O(n25430) );
  AO12S U21286 ( .B1(n25444), .B2(n25477), .A1(n25401), .O(n15293) );
  MUX2S U21287 ( .A(n28534), .B(n25475), .S(gray_img[1886]), .O(n25401) );
  AO12S U21288 ( .B1(n25444), .B2(n25460), .A1(n25391), .O(n15294) );
  MUX2S U21289 ( .A(n27447), .B(n25458), .S(gray_img[1878]), .O(n25391) );
  AO12S U21290 ( .B1(n25444), .B2(n25631), .A1(n25424), .O(n15295) );
  MUX2S U21291 ( .A(n28534), .B(n25629), .S(gray_img[1870]), .O(n25424) );
  ND2S U21292 ( .I1(n20022), .I2(n20021), .O(n15296) );
  MUX2S U21293 ( .A(n29587), .B(n20504), .S(gray_img[1862]), .O(n20021) );
  ND2S U21294 ( .I1(n20409), .I2(n20408), .O(n15297) );
  MUX2S U21295 ( .A(n29566), .B(n20740), .S(gray_img[1854]), .O(n20408) );
  ND2S U21296 ( .I1(n20372), .I2(n20371), .O(n15298) );
  MUX2S U21297 ( .A(n29597), .B(n20862), .S(gray_img[1846]), .O(n20372) );
  ND2S U21298 ( .I1(n20012), .I2(n20011), .O(n15299) );
  ND2S U21299 ( .I1(n20000), .I2(n19999), .O(n15300) );
  ND2S U21300 ( .I1(n20298), .I2(n20297), .O(n15301) );
  MUX2S U21301 ( .A(n29587), .B(n20296), .S(gray_img[1822]), .O(n20298) );
  ND2S U21302 ( .I1(n20351), .I2(n20350), .O(n15302) );
  MUX2S U21303 ( .A(n29597), .B(n20354), .S(gray_img[1814]), .O(n20351) );
  ND2S U21304 ( .I1(n20321), .I2(n20320), .O(n15303) );
  MUX2S U21305 ( .A(n30056), .B(n20319), .S(gray_img[1806]), .O(n20320) );
  MUX2S U21306 ( .A(n29597), .B(n20376), .S(gray_img[1798]), .O(n20378) );
  ND2S U21307 ( .I1(n20439), .I2(n20438), .O(n15305) );
  MUX2S U21308 ( .A(n29597), .B(n20547), .S(gray_img[1790]), .O(n20438) );
  ND2S U21309 ( .I1(n20448), .I2(n20447), .O(n15306) );
  MUX2S U21310 ( .A(n29566), .B(n20541), .S(gray_img[1782]), .O(n20447) );
  ND2S U21311 ( .I1(n20451), .I2(n20450), .O(n15307) );
  MUX2S U21312 ( .A(n30044), .B(n20449), .S(gray_img[1774]), .O(n20450) );
  AO12S U21313 ( .B1(n25444), .B2(n25778), .A1(n25435), .O(n15308) );
  MUX2S U21314 ( .A(n28534), .B(n25776), .S(gray_img[1766]), .O(n25435) );
  AO12S U21315 ( .B1(n25389), .B2(n25510), .A1(n25384), .O(n15309) );
  MUX2S U21316 ( .A(n27447), .B(n25508), .S(gray_img[1758]), .O(n25384) );
  AO12S U21317 ( .B1(n25444), .B2(n25498), .A1(n25429), .O(n15310) );
  AO12S U21318 ( .B1(n25389), .B2(n25649), .A1(n25387), .O(n15311) );
  MUX2S U21319 ( .A(n27447), .B(n25647), .S(gray_img[1742]), .O(n25387) );
  MUX2S U21320 ( .A(n29566), .B(n19955), .S(gray_img[1734]), .O(n18991) );
  ND2S U21321 ( .I1(n20405), .I2(n20404), .O(n15313) );
  MUX2S U21322 ( .A(n30044), .B(n20737), .S(gray_img[1726]), .O(n20404) );
  ND2S U21323 ( .I1(n20401), .I2(n20400), .O(n15314) );
  MUX2S U21324 ( .A(n30050), .B(n20846), .S(gray_img[1718]), .O(n20401) );
  ND2S U21325 ( .I1(n20008), .I2(n20007), .O(n15315) );
  MUX2S U21326 ( .A(n30056), .B(n20827), .S(gray_img[1710]), .O(n20008) );
  ND2S U21327 ( .I1(n20282), .I2(n20281), .O(n15316) );
  MUX2S U21328 ( .A(n30056), .B(n20787), .S(gray_img[1702]), .O(n20282) );
  ND2S U21329 ( .I1(n20383), .I2(n20382), .O(n15317) );
  MUX2S U21330 ( .A(n30044), .B(n20599), .S(gray_img[1694]), .O(n20383) );
  ND2S U21331 ( .I1(n19996), .I2(n19995), .O(n15318) );
  MUX2S U21332 ( .A(n29587), .B(n20605), .S(gray_img[1686]), .O(n19996) );
  ND2S U21333 ( .I1(n20315), .I2(n20314), .O(n15319) );
  MUX2S U21334 ( .A(n29566), .B(n20531), .S(gray_img[1678]), .O(n20314) );
  ND2S U21335 ( .I1(n20300), .I2(n20299), .O(n15320) );
  MUX2S U21336 ( .A(n29587), .B(n20583), .S(gray_img[1670]), .O(n20300) );
  ND2S U21337 ( .I1(n20462), .I2(n20461), .O(n15321) );
  ND2S U21338 ( .I1(n18563), .I2(n18562), .O(n15322) );
  MUX2S U21339 ( .A(n15904), .B(n20525), .S(gray_img[1654]), .O(n18562) );
  AO12S U21340 ( .B1(n25444), .B2(n25899), .A1(n25443), .O(n15324) );
  MUX2S U21341 ( .A(n27447), .B(n25897), .S(gray_img[1638]), .O(n25443) );
  AO12S U21342 ( .B1(n25389), .B2(n25576), .A1(n25382), .O(n15325) );
  MUX2S U21343 ( .A(n27447), .B(n25574), .S(gray_img[1630]), .O(n25382) );
  AO12S U21344 ( .B1(n25448), .B2(n25494), .A1(n25417), .O(n15326) );
  MUX2S U21345 ( .A(n28534), .B(n25492), .S(gray_img[1622]), .O(n25417) );
  AO12S U21346 ( .B1(n25448), .B2(n25653), .A1(n25380), .O(n15327) );
  MUX2S U21347 ( .A(n28534), .B(n25651), .S(gray_img[1614]), .O(n25380) );
  MUX2S U21348 ( .A(n29587), .B(n20528), .S(gray_img[1606]), .O(n18993) );
  ND2S U21349 ( .I1(n20411), .I2(n20410), .O(n15329) );
  MUX2S U21350 ( .A(n30056), .B(n20731), .S(gray_img[1598]), .O(n20410) );
  ND2S U21351 ( .I1(n20388), .I2(n20387), .O(n15330) );
  MUX2S U21352 ( .A(n20830), .B(n20839), .S(gray_img[1590]), .O(n20388) );
  ND2S U21353 ( .I1(n20397), .I2(n20396), .O(n15331) );
  MUX2S U21354 ( .A(n30050), .B(n20395), .S(gray_img[1582]), .O(n20397) );
  ND2S U21355 ( .I1(n19998), .I2(n19997), .O(n15332) );
  MUX2S U21356 ( .A(n30056), .B(n20824), .S(gray_img[1574]), .O(n19998) );
  MUX2S U21357 ( .A(n29597), .B(n20596), .S(gray_img[1566]), .O(n18615) );
  ND2S U21358 ( .I1(n20004), .I2(n20003), .O(n15334) );
  MUX2S U21359 ( .A(n29587), .B(n20602), .S(gray_img[1558]), .O(n20004) );
  MUX2S U21360 ( .A(n29566), .B(n20550), .S(gray_img[1550]), .O(n18716) );
  ND2S U21361 ( .I1(n20880), .I2(n20879), .O(n15336) );
  MUX2S U21362 ( .A(n29597), .B(n20881), .S(gray_img[1542]), .O(n20880) );
  ND2S U21363 ( .I1(n20407), .I2(n20406), .O(n15337) );
  MUX2S U21364 ( .A(n30056), .B(n20556), .S(gray_img[1534]), .O(n20406) );
  ND2S U21365 ( .I1(n20476), .I2(n20475), .O(n15338) );
  MUX2S U21366 ( .A(n30050), .B(n20440), .S(gray_img[1518]), .O(n20441) );
  AO12S U21367 ( .B1(n25448), .B2(n27971), .A1(n25447), .O(n15340) );
  MUX2S U21368 ( .A(n28534), .B(n27969), .S(gray_img[1510]), .O(n25447) );
  AO12S U21369 ( .B1(n25448), .B2(n28355), .A1(n25425), .O(n15341) );
  MUX2S U21370 ( .A(n15889), .B(n28353), .S(gray_img[1502]), .O(n25425) );
  AO12S U21371 ( .B1(n25448), .B2(n28342), .A1(n25408), .O(n15342) );
  AO12S U21372 ( .B1(n25448), .B2(n28560), .A1(n25406), .O(n15343) );
  ND2S U21373 ( .I1(n20415), .I2(n20414), .O(n15344) );
  MUX2S U21374 ( .A(n15904), .B(n20684), .S(gray_img[1478]), .O(n20414) );
  ND2S U21375 ( .I1(n20306), .I2(n20305), .O(n15345) );
  ND2S U21376 ( .I1(n20286), .I2(n20285), .O(n15346) );
  MUX2S U21377 ( .A(n30044), .B(n20821), .S(gray_img[1462]), .O(n20286) );
  ND2S U21378 ( .I1(n20010), .I2(n20009), .O(n15347) );
  MUX2S U21379 ( .A(n15904), .B(n20814), .S(gray_img[1454]), .O(n20010) );
  ND2S U21380 ( .I1(n20290), .I2(n20289), .O(n15348) );
  MUX2S U21381 ( .A(n30005), .B(n20811), .S(gray_img[1446]), .O(n20290) );
  ND2S U21382 ( .I1(n20295), .I2(n20294), .O(n15349) );
  MUX2S U21383 ( .A(n30044), .B(n20293), .S(gray_img[1438]), .O(n20295) );
  ND2S U21384 ( .I1(n18892), .I2(n18891), .O(n15350) );
  MUX2S U21385 ( .A(n20842), .B(n20193), .S(gray_img[1430]), .O(n18892) );
  ND2S U21386 ( .I1(n20018), .I2(n20017), .O(n15351) );
  MUX2S U21387 ( .A(n15904), .B(n20035), .S(gray_img[1422]), .O(n20017) );
  ND2S U21388 ( .I1(n20361), .I2(n20360), .O(n15352) );
  MUX2S U21389 ( .A(n20830), .B(n20359), .S(gray_img[1414]), .O(n20361) );
  MUX2S U21390 ( .A(n30050), .B(n20571), .S(gray_img[1406]), .O(n18755) );
  MUX2S U21391 ( .A(n30050), .B(n20517), .S(gray_img[1398]), .O(n20420) );
  ND2S U21392 ( .I1(n20456), .I2(n20455), .O(n15355) );
  MUX2S U21393 ( .A(n30050), .B(n20722), .S(gray_img[1390]), .O(n20455) );
  ND2S U21394 ( .I1(n15889), .I2(n27997), .O(n25440) );
  AO12S U21395 ( .B1(n25448), .B2(n28359), .A1(n25392), .O(n15357) );
  AO12S U21396 ( .B1(n25448), .B2(n28596), .A1(n25410), .O(n15358) );
  MUX2S U21397 ( .A(n15889), .B(n28594), .S(gray_img[1366]), .O(n25410) );
  AO12S U21398 ( .B1(n25444), .B2(n28536), .A1(n25407), .O(n15359) );
  ND2S U21399 ( .I1(n18990), .I2(n18989), .O(n15360) );
  MUX2S U21400 ( .A(n15904), .B(n20734), .S(gray_img[1350]), .O(n18989) );
  ND2S U21401 ( .I1(n20304), .I2(n20303), .O(n15361) );
  ND2S U21402 ( .I1(n20280), .I2(n20279), .O(n15362) );
  MUX2S U21403 ( .A(n30050), .B(n20833), .S(gray_img[1334]), .O(n20280) );
  ND2S U21404 ( .I1(n20002), .I2(n20001), .O(n15363) );
  MUX2S U21405 ( .A(n29566), .B(n20836), .S(gray_img[1326]), .O(n20002) );
  ND2S U21406 ( .I1(n20284), .I2(n20283), .O(n15364) );
  MUX2S U21407 ( .A(n29566), .B(n20843), .S(gray_img[1318]), .O(n20284) );
  ND2S U21408 ( .I1(n20014), .I2(n20013), .O(n15365) );
  ND2S U21409 ( .I1(n20364), .I2(n20363), .O(n15366) );
  MUX2S U21410 ( .A(n30056), .B(n20362), .S(gray_img[1302]), .O(n20364) );
  ND2S U21411 ( .I1(n20429), .I2(n20428), .O(n15367) );
  MUX2S U21412 ( .A(n20842), .B(n20427), .S(gray_img[1294]), .O(n20428) );
  ND2S U21413 ( .I1(n20394), .I2(n20393), .O(n15368) );
  MUX2S U21414 ( .A(n15904), .B(n20392), .S(gray_img[1286]), .O(n20394) );
  ND2S U21415 ( .I1(n20308), .I2(n20307), .O(n15369) );
  ND2S U21416 ( .I1(n18588), .I2(n18587), .O(n15370) );
  MUX2S U21417 ( .A(n20808), .B(n20725), .S(gray_img[1270]), .O(n18587) );
  MUX2S U21418 ( .A(n30056), .B(n20719), .S(gray_img[1262]), .O(n18966) );
  AO12S U21419 ( .B1(n25444), .B2(n28031), .A1(n25431), .O(n15372) );
  MUX2S U21420 ( .A(n15889), .B(n28029), .S(gray_img[1254]), .O(n25431) );
  AO12S U21421 ( .B1(n25448), .B2(n28288), .A1(n25428), .O(n15373) );
  AO12S U21422 ( .B1(n25389), .B2(n28271), .A1(n25388), .O(n15374) );
  MUX2S U21423 ( .A(n15889), .B(n28269), .S(gray_img[1238]), .O(n25388) );
  AO12S U21424 ( .B1(n25448), .B2(n28475), .A1(n25416), .O(n15375) );
  MUX2S U21425 ( .A(n29587), .B(n20702), .S(gray_img[1222]), .O(n20433) );
  ND2S U21426 ( .I1(n20020), .I2(n20019), .O(n15377) );
  MUX2S U21427 ( .A(n30044), .B(n20757), .S(gray_img[1214]), .O(n20019) );
  ND2S U21428 ( .I1(n20288), .I2(n20287), .O(n15378) );
  MUX2S U21429 ( .A(n30044), .B(n20857), .S(gray_img[1206]), .O(n20288) );
  ND2S U21430 ( .I1(n20437), .I2(n20436), .O(n15379) );
  MUX2S U21431 ( .A(n29566), .B(n20435), .S(gray_img[1198]), .O(n20436) );
  MUX2S U21432 ( .A(n29566), .B(n20379), .S(gray_img[1190]), .O(n20381) );
  MUX2S U21433 ( .A(n29597), .B(n20159), .S(gray_img[1182]), .O(n18620) );
  ND2S U21434 ( .I1(n20318), .I2(n20317), .O(n15382) );
  MUX2S U21435 ( .A(n30005), .B(n20316), .S(gray_img[1174]), .O(n20317) );
  ND2S U21436 ( .I1(n20016), .I2(n20015), .O(n15383) );
  MUX2S U21437 ( .A(n30044), .B(n20553), .S(gray_img[1166]), .O(n20015) );
  ND2S U21438 ( .I1(n20024), .I2(n20023), .O(n15384) );
  MUX2S U21439 ( .A(n30056), .B(n20240), .S(gray_img[1158]), .O(n20023) );
  MUX2S U21440 ( .A(n30056), .B(n20716), .S(gray_img[1150]), .O(n20470) );
  ND2S U21441 ( .I1(n18591), .I2(n18590), .O(n15386) );
  MUX2S U21442 ( .A(n20808), .B(n20124), .S(gray_img[1142]), .O(n18590) );
  MUX2S U21443 ( .A(n30044), .B(n20728), .S(gray_img[1134]), .O(n18963) );
  AO12S U21444 ( .B1(n25448), .B2(n28092), .A1(n25445), .O(n15388) );
  MUX2S U21445 ( .A(n28534), .B(n28090), .S(gray_img[1126]), .O(n25445) );
  AO12S U21446 ( .B1(n25448), .B2(n28284), .A1(n25419), .O(n15389) );
  AO12S U21447 ( .B1(n25444), .B2(n28423), .A1(n25400), .O(n15390) );
  AO12S U21448 ( .B1(n25448), .B2(n28480), .A1(n25394), .O(n15391) );
  MUX2S U21449 ( .A(n15889), .B(n28478), .S(gray_img[1102]), .O(n25394) );
  MUX2S U21450 ( .A(n30050), .B(n20743), .S(gray_img[1094]), .O(n20443) );
  ND2S U21451 ( .I1(n20302), .I2(n20301), .O(n15393) );
  MUX2S U21452 ( .A(n30056), .B(n20760), .S(gray_img[1086]), .O(n20301) );
  ND2S U21453 ( .I1(n20292), .I2(n20291), .O(n15394) );
  MUX2S U21454 ( .A(n30044), .B(n20854), .S(gray_img[1078]), .O(n20292) );
  ND2S U21455 ( .I1(n20446), .I2(n20445), .O(n15395) );
  MUX2S U21456 ( .A(n29597), .B(n20611), .S(gray_img[1070]), .O(n20445) );
  MUX2S U21457 ( .A(n29587), .B(n20368), .S(gray_img[1062]), .O(n20370) );
  MUX2S U21458 ( .A(n29597), .B(n20184), .S(gray_img[1054]), .O(n18624) );
  ND2S U21459 ( .I1(n19779), .I2(n19778), .O(n15398) );
  MUX2S U21460 ( .A(n29587), .B(n20255), .S(gray_img[1046]), .O(n19778) );
  MUX2S U21461 ( .A(n29566), .B(n20235), .S(gray_img[1038]), .O(n19416) );
  ND2S U21462 ( .I1(n20313), .I2(n20312), .O(n15400) );
  MUX2S U21463 ( .A(n29587), .B(n20311), .S(gray_img[1030]), .O(n20312) );
  ND2S U21464 ( .I1(n18673), .I2(n18672), .O(n15401) );
  MUX2S U21465 ( .A(n30005), .B(n20099), .S(gray_img[1022]), .O(n18672) );
  ND2S U21466 ( .I1(n18565), .I2(n18564), .O(n15402) );
  MUX2S U21467 ( .A(n30005), .B(n20562), .S(gray_img[1014]), .O(n18564) );
  MUX2S U21468 ( .A(n20830), .B(n20384), .S(gray_img[1006]), .O(n20386) );
  AO12S U21469 ( .B1(n25444), .B2(n27829), .A1(n25436), .O(n15404) );
  AO12S U21470 ( .B1(n25444), .B2(n27081), .A1(n25397), .O(n15405) );
  MUX2S U21471 ( .A(n15889), .B(n27079), .S(gray_img[990]), .O(n25397) );
  AO12S U21472 ( .B1(n25448), .B2(n27065), .A1(n25393), .O(n15406) );
  MUX2S U21473 ( .A(n15889), .B(n27063), .S(gray_img[982]), .O(n25393) );
  AO12S U21474 ( .B1(n25444), .B2(n27261), .A1(n25409), .O(n15407) );
  MUX2S U21475 ( .A(n29587), .B(n20580), .S(gray_img[966]), .O(n18933) );
  ND2S U21476 ( .I1(n20454), .I2(n20453), .O(n15409) );
  MUX2S U21477 ( .A(n30005), .B(n20452), .S(gray_img[894]), .O(n20453) );
  ND2S U21478 ( .I1(n20310), .I2(n20309), .O(n15410) );
  MUX2S U21479 ( .A(n30005), .B(n20559), .S(gray_img[886]), .O(n20309) );
  ND2S U21480 ( .I1(n18914), .I2(n18913), .O(n15411) );
  MUX2S U21481 ( .A(n30005), .B(n20212), .S(gray_img[878]), .O(n18914) );
  AO12S U21482 ( .B1(n25444), .B2(n26224), .A1(n25432), .O(n15412) );
  MUX2S U21483 ( .A(n28534), .B(n26222), .S(gray_img[870]), .O(n25432) );
  AO12S U21484 ( .B1(n25448), .B2(n30065), .A1(n25413), .O(n15413) );
  AO12S U21485 ( .B1(n25444), .B2(n27069), .A1(n25421), .O(n15414) );
  AO12S U21486 ( .B1(n25448), .B2(n27190), .A1(n25390), .O(n15415) );
  ND2S U21487 ( .I1(n20458), .I2(n20457), .O(n15416) );
  MUX2S U21488 ( .A(n20634), .B(n30005), .S(n22971), .O(n20457) );
  ND2S U21489 ( .I1(n20460), .I2(n20459), .O(n15417) );
  MUX2S U21490 ( .A(n30005), .B(n20568), .S(gray_img[766]), .O(n20459) );
  ND2S U21491 ( .I1(n18559), .I2(n18558), .O(n15418) );
  MUX2S U21492 ( .A(n15904), .B(n20054), .S(gray_img[758]), .O(n18558) );
  ND2S U21493 ( .I1(n20367), .I2(n20366), .O(n15419) );
  MUX2S U21494 ( .A(n30005), .B(n20365), .S(gray_img[750]), .O(n20367) );
  AO12S U21495 ( .B1(n25448), .B2(n26155), .A1(n25437), .O(n15420) );
  AO12S U21496 ( .B1(n25444), .B2(n26996), .A1(n25415), .O(n15421) );
  MUX2S U21497 ( .A(n15889), .B(n26994), .S(gray_img[734]), .O(n25415) );
  AO12S U21498 ( .B1(n25448), .B2(n27009), .A1(n25396), .O(n15422) );
  AO12S U21499 ( .B1(n25448), .B2(n27243), .A1(n25420), .O(n15423) );
  ND2S U21500 ( .I1(n19873), .I2(n19872), .O(n15424) );
  MUX2S U21501 ( .A(n29587), .B(n20623), .S(gray_img[710]), .O(n19872) );
  ND2S U21502 ( .I1(n20467), .I2(n20466), .O(n15425) );
  MUX2S U21503 ( .A(n25928), .B(n20565), .S(gray_img[638]), .O(n20466) );
  ND2S U21504 ( .I1(n20469), .I2(n20468), .O(n15426) );
  MUX2S U21505 ( .A(n30050), .B(n20534), .S(gray_img[630]), .O(n20468) );
  ND2S U21506 ( .I1(n19841), .I2(n19840), .O(n15427) );
  MUX2S U21507 ( .A(n15904), .B(n20274), .S(gray_img[622]), .O(n19840) );
  AO12S U21508 ( .B1(n25448), .B2(n26160), .A1(n25433), .O(n15428) );
  AO12S U21509 ( .B1(n25444), .B2(n27105), .A1(n25418), .O(n15429) );
  AO12S U21510 ( .B1(n25389), .B2(n27013), .A1(n25385), .O(n15430) );
  AO12S U21511 ( .B1(n25444), .B2(n27133), .A1(n25398), .O(n15431) );
  MUX2S U21512 ( .A(n29566), .B(n20591), .S(gray_img[582]), .O(n20399) );
  MUX2S U21513 ( .A(n30050), .B(n20472), .S(gray_img[510]), .O(n20473) );
  ND2S U21514 ( .I1(n20479), .I2(n20478), .O(n15434) );
  MUX2S U21515 ( .A(n30056), .B(n20477), .S(gray_img[502]), .O(n20478) );
  ND2S U21516 ( .I1(n20482), .I2(n20481), .O(n15435) );
  MUX2S U21517 ( .A(n29566), .B(n20480), .S(gray_img[494]), .O(n20481) );
  AO12S U21518 ( .B1(n25448), .B2(n27774), .A1(n25446), .O(n15436) );
  MUX2S U21519 ( .A(n27447), .B(n27772), .S(gray_img[486]), .O(n25446) );
  AO12S U21520 ( .B1(n25389), .B2(n27352), .A1(n25383), .O(n15437) );
  MUX2S U21521 ( .A(n27447), .B(n27350), .S(gray_img[478]), .O(n25383) );
  AO12S U21522 ( .B1(n25444), .B2(n26747), .A1(n25379), .O(n15438) );
  MUX2S U21523 ( .A(n28534), .B(n26745), .S(gray_img[470]), .O(n25379) );
  AO12S U21524 ( .B1(n25448), .B2(n26942), .A1(n25427), .O(n15439) );
  ND2S U21525 ( .I1(n20485), .I2(n20484), .O(n15440) );
  MUX2S U21526 ( .A(n30005), .B(n20483), .S(gray_img[454]), .O(n20484) );
  ND2S U21527 ( .I1(n20488), .I2(n20487), .O(n15441) );
  MUX2S U21528 ( .A(n30056), .B(n20486), .S(gray_img[382]), .O(n20487) );
  MUX2S U21529 ( .A(n30050), .B(n20522), .S(gray_img[374]), .O(n20489) );
  ND2S U21530 ( .I1(n20493), .I2(n20492), .O(n15443) );
  MUX2S U21531 ( .A(n29566), .B(n20491), .S(gray_img[366]), .O(n20492) );
  AO12S U21532 ( .B1(n25444), .B2(n27449), .A1(n25438), .O(n15444) );
  MUX2S U21533 ( .A(n28534), .B(n27446), .S(gray_img[358]), .O(n25438) );
  AO12S U21534 ( .B1(n25448), .B2(n26759), .A1(n25426), .O(n15445) );
  AO12S U21535 ( .B1(n25448), .B2(n26743), .A1(n25402), .O(n15446) );
  MUX2S U21536 ( .A(n28534), .B(n26741), .S(gray_img[342]), .O(n25402) );
  AO12S U21537 ( .B1(n25448), .B2(n26861), .A1(n25423), .O(n15447) );
  MUX2S U21538 ( .A(n27447), .B(n26859), .S(gray_img[334]), .O(n25423) );
  ND2S U21539 ( .I1(n18935), .I2(n18934), .O(n15448) );
  MUX2S U21540 ( .A(n30005), .B(n20147), .S(gray_img[326]), .O(n18935) );
  MUX2S U21541 ( .A(n29566), .B(n20496), .S(gray_img[254]), .O(n20497) );
  ND2S U21542 ( .I1(n19735), .I2(n19734), .O(n15450) );
  MUX2S U21543 ( .A(n30056), .B(n20260), .S(gray_img[246]), .O(n19734) );
  MUX2S U21544 ( .A(n20620), .B(n20830), .S(n27405), .O(n20494) );
  AO12S U21545 ( .B1(n25444), .B2(n27390), .A1(n25442), .O(n15452) );
  MUX2S U21546 ( .A(n27447), .B(n27388), .S(gray_img[230]), .O(n25442) );
  AO12S U21547 ( .B1(n25389), .B2(n26726), .A1(n25386), .O(n15453) );
  AO12S U21548 ( .B1(n25448), .B2(n26841), .A1(n25399), .O(n15454) );
  AO12S U21549 ( .B1(n25448), .B2(n26883), .A1(n25412), .O(n15455) );
  MUX2S U21550 ( .A(n15889), .B(n26881), .S(gray_img[206]), .O(n25412) );
  ND2S U21551 ( .I1(n19893), .I2(n19892), .O(n15456) );
  MUX2S U21552 ( .A(n15904), .B(n20631), .S(gray_img[198]), .O(n19892) );
  MUX2S U21553 ( .A(n30056), .B(n20082), .S(gray_img[126]), .O(n18646) );
  ND2S U21554 ( .I1(n20501), .I2(n20500), .O(n15458) );
  MUX2S U21555 ( .A(n30044), .B(n20499), .S(gray_img[118]), .O(n20500) );
  ND2S U21556 ( .I1(n20503), .I2(n20502), .O(n15459) );
  MUX2S U21557 ( .A(n20617), .B(n20830), .S(n27401), .O(n20502) );
  AO12S U21558 ( .B1(n25444), .B2(n27545), .A1(n25434), .O(n15460) );
  MUX2S U21559 ( .A(n28534), .B(n27543), .S(gray_img[102]), .O(n25434) );
  AO12S U21560 ( .B1(n25444), .B2(n26709), .A1(n25395), .O(n15461) );
  MUX2S U21561 ( .A(n15889), .B(n26707), .S(gray_img[94]), .O(n25395) );
  AO12S U21562 ( .B1(n25448), .B2(n26722), .A1(n25411), .O(n15462) );
  AO12S U21563 ( .B1(n25444), .B2(n26879), .A1(n25422), .O(n15463) );
  MUX2S U21564 ( .A(n28534), .B(n26877), .S(gray_img[78]), .O(n25422) );
  ND2S U21565 ( .I1(n19908), .I2(n19907), .O(n15464) );
  MUX2S U21566 ( .A(n15904), .B(n20628), .S(gray_img[70]), .O(n19907) );
  ND2S U21567 ( .I1(n21336), .I2(n21335), .O(n15809) );
  ND2S U21568 ( .I1(n30120), .I2(n23473), .O(n23476) );
  MUX2S U21569 ( .A(template_in_reg[7]), .B(template_reg[47]), .S(n30141), .O(
        n15685) );
  MUX2S U21570 ( .A(template_in_reg[6]), .B(template_reg[46]), .S(n30141), .O(
        n15686) );
  MUX2S U21571 ( .A(template_in_reg[5]), .B(template_reg[45]), .S(n30141), .O(
        n15687) );
  MUX2S U21572 ( .A(template_in_reg[4]), .B(template_reg[44]), .S(n30141), .O(
        n15688) );
  MUX2S U21573 ( .A(template_in_reg[3]), .B(template_reg[43]), .S(n30141), .O(
        n15689) );
  MUX2S U21574 ( .A(template_in_reg[2]), .B(template_reg[42]), .S(n30141), .O(
        n15690) );
  MUX2S U21575 ( .A(template_in_reg[1]), .B(template_reg[41]), .S(n30141), .O(
        n15691) );
  MUX2S U21576 ( .A(template_in_reg[0]), .B(template_reg[40]), .S(n30141), .O(
        n15692) );
  MUX2S U21577 ( .A(template_in_reg[7]), .B(template_reg[39]), .S(n30140), .O(
        n15693) );
  MUX2S U21578 ( .A(template_in_reg[6]), .B(template_reg[38]), .S(n30140), .O(
        n15694) );
  MUX2S U21579 ( .A(template_in_reg[5]), .B(template_reg[37]), .S(n30140), .O(
        n15695) );
  MUX2S U21580 ( .A(template_in_reg[4]), .B(template_reg[36]), .S(n30140), .O(
        n15696) );
  MUX2S U21581 ( .A(template_in_reg[3]), .B(template_reg[35]), .S(n30140), .O(
        n15697) );
  MUX2S U21582 ( .A(template_in_reg[2]), .B(template_reg[34]), .S(n30140), .O(
        n15698) );
  MUX2S U21583 ( .A(template_in_reg[1]), .B(template_reg[33]), .S(n30140), .O(
        n15699) );
  MUX2S U21584 ( .A(template_in_reg[0]), .B(template_reg[32]), .S(n30140), .O(
        n15700) );
  MUX2S U21585 ( .A(template_in_reg[7]), .B(template_reg[31]), .S(n30142), .O(
        n15701) );
  MUX2S U21586 ( .A(template_in_reg[6]), .B(template_reg[30]), .S(n30142), .O(
        n15702) );
  MUX2S U21587 ( .A(template_in_reg[5]), .B(template_reg[29]), .S(n30142), .O(
        n15703) );
  MUX2S U21588 ( .A(template_in_reg[4]), .B(template_reg[28]), .S(n30142), .O(
        n15704) );
  MUX2S U21589 ( .A(template_in_reg[3]), .B(template_reg[27]), .S(n30142), .O(
        n15705) );
  MUX2S U21590 ( .A(template_in_reg[2]), .B(template_reg[26]), .S(n30142), .O(
        n15706) );
  MUX2S U21591 ( .A(template_in_reg[1]), .B(template_reg[25]), .S(n30142), .O(
        n15707) );
  MUX2S U21592 ( .A(template_in_reg[0]), .B(template_reg[24]), .S(n30142), .O(
        n15708) );
  BUF1CK U21593 ( .I(medfilt_state[1]), .O(n30453) );
  OR2 U21594 ( .I1(n16208), .I2(n16213), .O(n15941) );
  BUF2 U21595 ( .I(n16380), .O(n17807) );
  OR2 U21596 ( .I1(n16164), .I2(n16173), .O(n15942) );
  AN2 U21597 ( .I1(n16974), .I2(n16973), .O(n15943) );
  OR2 U21598 ( .I1(n16211), .I2(n16207), .O(n15944) );
  AN2 U21599 ( .I1(n17822), .I2(n17821), .O(n15945) );
  NR2T U21600 ( .I1(n16212), .I2(n16196), .O(n16188) );
  INV3 U21601 ( .I(n15998), .O(n17796) );
  OR2 U21602 ( .I1(n16168), .I2(n16209), .O(n15946) );
  BUF2 U21603 ( .I(n16121), .O(n17703) );
  OR2 U21604 ( .I1(n16198), .I2(n16207), .O(n15947) );
  INV2 U21605 ( .I(n15999), .O(n17752) );
  NR2T U21606 ( .I1(n16207), .I2(n16168), .O(n15948) );
  NR2T U21607 ( .I1(n16205), .I2(n16209), .O(n16116) );
  INV3 U21608 ( .I(n16477), .O(n17605) );
  NR2T U21609 ( .I1(n16207), .I2(n16205), .O(n15949) );
  NR2T U21610 ( .I1(n16213), .I2(n16212), .O(n15950) );
  NR2T U21611 ( .I1(n16207), .I2(n16212), .O(n15951) );
  NR2P U21612 ( .I1(n24755), .I2(n24798), .O(n24855) );
  FA1 U21613 ( .A(n17912), .B(n17911), .CI(n17910), .CO(n17916), .S(n17908) );
  FA1S U21614 ( .A(n17906), .B(n17905), .CI(n17904), .CO(n17910), .S(n17894)
         );
  XOR2HS U21615 ( .I1(cnt_cro_3b3[0]), .I2(cnt_cro_y[0]), .O(n16157) );
  ND2P U21616 ( .I1(n16148), .I2(n16147), .O(n16151) );
  OR2S U21617 ( .I1(n28077), .I2(n28079), .O(n15963) );
  NR2 U21618 ( .I1(n29680), .I2(n16045), .O(n26849) );
  OR2S U21619 ( .I1(n28542), .I2(n28540), .O(n15976) );
  OR2S U21620 ( .I1(n27808), .I2(n27806), .O(n15977) );
  OA112S U21621 ( .C1(n24653), .C2(n24380), .A1(n24356), .B1(n24355), .O(
        n15985) );
  OR2 U21622 ( .I1(n24513), .I2(n24241), .O(n15986) );
  AN2 U21623 ( .I1(n24252), .I2(n24253), .O(n15987) );
  AN2 U21624 ( .I1(n24143), .I2(n24353), .O(n15988) );
  AN2S U21625 ( .I1(n24652), .I2(n24353), .O(n15989) );
  AOI12HS U21626 ( .B1(n24951), .B2(n17590), .A1(n17589), .O(n15990) );
  AOI12HS U21627 ( .B1(n24951), .B2(n17363), .A1(n17362), .O(n15991) );
  AOI12HS U21628 ( .B1(n24951), .B2(n16096), .A1(n16095), .O(n15992) );
  AOI12HS U21629 ( .B1(n24951), .B2(n16402), .A1(n16401), .O(n15993) );
  AOI12HS U21630 ( .B1(n24951), .B2(n16596), .A1(n16595), .O(n15994) );
  AOI12HS U21631 ( .B1(n24951), .B2(n16980), .A1(n16979), .O(n15995) );
  AOI12HS U21632 ( .B1(n24951), .B2(n16792), .A1(n16791), .O(n15996) );
  AOI12HS U21633 ( .B1(n24951), .B2(n16602), .A1(n16601), .O(n15997) );
  OR2 U21634 ( .I1(n16211), .I2(n16204), .O(n15998) );
  OR2 U21635 ( .I1(n16211), .I2(n16174), .O(n15999) );
  OR2 U21636 ( .I1(n16208), .I2(n16204), .O(n16379) );
  NR2 U21637 ( .I1(n16210), .I2(n16174), .O(n16500) );
  NR2T U21638 ( .I1(n16198), .I2(n16204), .O(n17805) );
  NR2 U21639 ( .I1(n16198), .I2(n16173), .O(n16296) );
  NR2T U21640 ( .I1(n16208), .I2(n16173), .O(n16000) );
  OR2 U21641 ( .I1(n16211), .I2(n16173), .O(n16495) );
  BUF2 U21642 ( .I(n17798), .O(n17717) );
  BUF2 U21643 ( .I(n17798), .O(n17606) );
  NR2T U21644 ( .I1(n16198), .I2(n16213), .O(n16001) );
  OR2 U21645 ( .I1(n16208), .I2(n16203), .O(n16002) );
  OA112S U21646 ( .C1(n26846), .C2(n16068), .A1(n16067), .B1(n16066), .O(
        n16004) );
  OA112S U21647 ( .C1(n26846), .C2(n16060), .A1(n16059), .B1(n16058), .O(
        n16005) );
  NR2P U21648 ( .I1(n16113), .I2(n16112), .O(n16114) );
  INV2 U21649 ( .I(n15941), .O(n17137) );
  AOI22S U21650 ( .A1(n17744), .A2(gray_img[565]), .B1(n16137), .B2(
        gray_img[813]), .O(n17072) );
  INV1S U21651 ( .I(n16280), .O(n17533) );
  AN4B1S U21652 ( .I1(n17127), .I2(n17126), .I3(n17125), .B1(n17124), .O(
        n17134) );
  AN4B1S U21653 ( .I1(n17074), .I2(n17073), .I3(n17072), .B1(n17071), .O(
        n17092) );
  INV1S U21654 ( .I(n16207), .O(n16122) );
  AN4B1S U21655 ( .I1(n16146), .I2(n16145), .I3(n16144), .B1(n16143), .O(
        n16180) );
  BUF2 U21656 ( .I(n16280), .O(n17806) );
  INV2 U21657 ( .I(n16668), .O(n17804) );
  INV3 U21658 ( .I(n15942), .O(n17751) );
  BUF2 U21659 ( .I(n16139), .O(n17709) );
  AOI12HS U21660 ( .B1(n24151), .B2(n24150), .A1(n24149), .O(n24154) );
  INV1S U21661 ( .I(gray_img[929]), .O(n23220) );
  ND3S U21662 ( .I1(n16978), .I2(n16977), .I3(n16976), .O(n16979) );
  INV1S U21663 ( .I(n24254), .O(n24228) );
  INV1S U21664 ( .I(gray_img[153]), .O(n27864) );
  INV1S U21665 ( .I(gray_img[817]), .O(n26098) );
  MAO222S U21666 ( .A1(gray_img[1665]), .B1(gray_img[1664]), .C1(n26588), .O(
        n26589) );
  MAO222S U21667 ( .A1(gray_img[1433]), .B1(gray_img[1432]), .C1(n29760), .O(
        n29761) );
  MAO222S U21668 ( .A1(gray_img[1073]), .B1(gray_img[1072]), .C1(n28866), .O(
        n28867) );
  INV1S U21669 ( .I(gray_img[1881]), .O(n23247) );
  ND3S U21670 ( .I1(n16600), .I2(n16599), .I3(n16598), .O(n16601) );
  ND3S U21671 ( .I1(n16400), .I2(n16399), .I3(n16398), .O(n16401) );
  AN4S U21672 ( .I1(n17739), .I2(n17738), .I3(n17737), .I4(n17736), .O(n17740)
         );
  OAI12HS U21673 ( .B1(n15989), .B2(n24007), .A1(n24006), .O(n24021) );
  NR2 U21674 ( .I1(n23847), .I2(n23854), .O(n23857) );
  ND3S U21675 ( .I1(n21477), .I2(n21476), .I3(n21475), .O(n21478) );
  ND3S U21676 ( .I1(n22816), .I2(n22815), .I3(n22814), .O(n22817) );
  MAO222S U21677 ( .A1(n28622), .B1(gray_img[674]), .C1(n28621), .O(n28623) );
  MAO222S U21678 ( .A1(gray_img[33]), .B1(gray_img[32]), .C1(n26943), .O(
        n26944) );
  NR2 U21679 ( .I1(n23641), .I2(n23687), .O(n23652) );
  NR2 U21680 ( .I1(n23649), .I2(n23687), .O(n23666) );
  INV1S U21681 ( .I(n17851), .O(n17854) );
  NR2 U21682 ( .I1(n16340), .I2(n16339), .O(n17690) );
  ND3S U21683 ( .I1(n22198), .I2(n22197), .I3(n22196), .O(n22199) );
  AOI12HS U21684 ( .B1(n24063), .B2(n24062), .A1(n24061), .O(n24064) );
  NR2 U21685 ( .I1(n23642), .I2(n23687), .O(n23645) );
  OAI12HS U21686 ( .B1(n23795), .B2(n23794), .A1(n23793), .O(n23796) );
  MAO222S U21687 ( .A1(n23142), .B1(gray_img[1843]), .C1(n23141), .O(n23143)
         );
  MAO222S U21688 ( .A1(n26550), .B1(gray_img[1555]), .C1(n26549), .O(n26551)
         );
  MAO222S U21689 ( .A1(n28964), .B1(gray_img[1322]), .C1(n28963), .O(n28965)
         );
  NR2 U21690 ( .I1(n23954), .I2(n23960), .O(n23958) );
  OAI12HS U21691 ( .B1(n23781), .B2(n24292), .A1(n23746), .O(n24547) );
  MOAI1S U21692 ( .A1(n17855), .A2(n17854), .B1(n17853), .B2(n17852), .O(
        n17933) );
  ND3S U21693 ( .I1(n17588), .I2(n17587), .I3(n17586), .O(n17589) );
  OA112S U21694 ( .C1(n22904), .C2(n26668), .A1(n21950), .B1(n21949), .O(
        n21951) );
  ND3S U21695 ( .I1(n21794), .I2(n21793), .I3(n21792), .O(n21795) );
  ND3S U21696 ( .I1(n22169), .I2(n22168), .I3(n22167), .O(n22170) );
  ND3S U21697 ( .I1(n22010), .I2(n22009), .I3(n22008), .O(n22011) );
  OA112S U21698 ( .C1(n26390), .C2(n22725), .A1(n22248), .B1(n22247), .O(
        n22250) );
  ND3S U21699 ( .I1(n21482), .I2(n21481), .I3(n21480), .O(n21484) );
  ND3S U21700 ( .I1(n21732), .I2(n21731), .I3(n21730), .O(n21748) );
  ND3S U21701 ( .I1(n21637), .I2(n21636), .I3(n21635), .O(n21638) );
  ND3S U21702 ( .I1(n22899), .I2(n22898), .I3(n22897), .O(n22916) );
  MAO222S U21703 ( .A1(n29391), .B1(gray_img[1923]), .C1(n29390), .O(n29392)
         );
  MOAI1S U21704 ( .A1(n24380), .A2(n24638), .B1(n24379), .B2(n24636), .O(
        n24362) );
  MOAI1S U21705 ( .A1(n24380), .A2(n24688), .B1(n24379), .B2(n24686), .O(
        n24371) );
  INV1S U21706 ( .I(mem_data_out_reg_shift_1[22]), .O(n24270) );
  ND3S U21707 ( .I1(n24693), .I2(n24172), .I3(n24354), .O(n24173) );
  INV1S U21708 ( .I(n22346), .O(n22802) );
  AOI12HS U21709 ( .B1(n24169), .B2(n24639), .A1(n24160), .O(n24199) );
  INV2 U21710 ( .I(n24427), .O(n24430) );
  INV1S U21711 ( .I(n21841), .O(n22566) );
  ND3S U21712 ( .I1(n22246), .I2(n22245), .I3(n22244), .O(n22253) );
  ND3S U21713 ( .I1(n21541), .I2(n21540), .I3(n21539), .O(n21542) );
  OA112S U21714 ( .C1(n22251), .C2(n29508), .A1(n21494), .B1(n21493), .O(
        n21497) );
  ND3S U21715 ( .I1(n21706), .I2(n21705), .I3(n21704), .O(n21707) );
  NR2 U21716 ( .I1(n23544), .I2(n23548), .O(n23531) );
  ND3S U21717 ( .I1(n21191), .I2(n21190), .I3(n21189), .O(n21192) );
  FA1S U21718 ( .A(n17983), .B(n17982), .CI(n17981), .CO(n17992), .S(n17989)
         );
  FA1S U21719 ( .A(n17986), .B(n17985), .CI(n17984), .CO(n17990), .S(n17966)
         );
  ND3S U21720 ( .I1(n21925), .I2(n21924), .I3(n21923), .O(n21926) );
  ND3S U21721 ( .I1(n22148), .I2(n22147), .I3(n22146), .O(n22149) );
  ND3S U21722 ( .I1(n22065), .I2(n22064), .I3(n22063), .O(n22096) );
  AO12 U21723 ( .B1(n24382), .B2(n24661), .A1(n24352), .O(n24418) );
  NR2 U21724 ( .I1(n24430), .I2(n24429), .O(n24608) );
  ND3S U21725 ( .I1(n22530), .I2(n22529), .I3(n22528), .O(n22531) );
  ND3S U21726 ( .I1(n22372), .I2(n22371), .I3(n22370), .O(n22373) );
  ND3S U21727 ( .I1(n21497), .I2(n21496), .I3(n21495), .O(n21498) );
  MOAI1S U21728 ( .A1(n27588), .A2(n27587), .B1(n27598), .B2(n27596), .O(
        n27589) );
  NR2 U21729 ( .I1(n24999), .I2(n25051), .O(n19913) );
  ND3S U21730 ( .I1(n24344), .I2(n24674), .I3(n24677), .O(n24407) );
  INV1S U21731 ( .I(n27375), .O(n27365) );
  AOI12HS U21732 ( .B1(n24331), .B2(n24285), .A1(n24284), .O(n24452) );
  ND3S U21733 ( .I1(n19402), .I2(n19401), .I3(n19400), .O(n19404) );
  NR2 U21734 ( .I1(n18884), .I2(n18822), .O(n25371) );
  INV1S U21735 ( .I(n28714), .O(n28717) );
  INV1S U21736 ( .I(n29593), .O(n29596) );
  INV1S U21737 ( .I(n24762), .O(n24859) );
  NR2 U21738 ( .I1(n18822), .I2(n25051), .O(n19719) );
  NR2 U21739 ( .I1(n25052), .I2(n25051), .O(n25339) );
  INV1S U21740 ( .I(cnt_cro_y[2]), .O(n25037) );
  INV2 U21741 ( .I(n19087), .O(n24069) );
  INV1S U21742 ( .I(in_valid), .O(n30387) );
  ND3S U21743 ( .I1(n21984), .I2(n21983), .I3(n21982), .O(n21985) );
  OA112S U21744 ( .C1(n24620), .C2(n24565), .A1(n24564), .B1(n24563), .O(
        n24867) );
  ND3S U21745 ( .I1(n21771), .I2(n21770), .I3(n21769), .O(n21772) );
  ND3S U21746 ( .I1(n22860), .I2(n22859), .I3(n22858), .O(n22958) );
  OR2 U21747 ( .I1(n29680), .I2(n26019), .O(n26077) );
  NR2 U21748 ( .I1(n29680), .I2(n23334), .O(n23492) );
  NR2 U21749 ( .I1(n29680), .I2(n23043), .O(n29043) );
  NR2 U21750 ( .I1(n29680), .I2(n27169), .O(n27251) );
  ND3S U21751 ( .I1(n25041), .I2(n25040), .I3(n30373), .O(n25034) );
  INV1S U21752 ( .I(image[2]), .O(n30416) );
  ND3S U21753 ( .I1(n18218), .I2(n18217), .I3(n18216), .O(n18223) );
  ND3S U21754 ( .I1(n28940), .I2(n28939), .I3(n28938), .O(n28941) );
  ND3S U21755 ( .I1(n18203), .I2(n18202), .I3(n18201), .O(n18212) );
  ND3S U21756 ( .I1(n18293), .I2(n18292), .I3(n18291), .O(n18294) );
  ND3S U21757 ( .I1(n18191), .I2(n18190), .I3(n18189), .O(n18200) );
  ND3S U21758 ( .I1(n18251), .I2(n18250), .I3(n18249), .O(n18260) );
  NR2 U21759 ( .I1(n29680), .I2(n29425), .O(n30098) );
  ND3S U21760 ( .I1(n19091), .I2(n24047), .I3(n18396), .O(n15806) );
  MOAI1S U21761 ( .A1(n30452), .A2(n30423), .B1(C551_DATA2_5), .B2(n30349), 
        .O(gray_scale_2_n[5]) );
  OAI112HS U21762 ( .C1(n18144), .C2(n30125), .A1(n18143), .B1(n18142), .O(
        n13623) );
  OAI112HS U21763 ( .C1(n18101), .C2(n29340), .A1(n18100), .B1(n18099), .O(
        n13953) );
  TIE1 U21764 ( .O(net76341) );
  OAI12HS U21765 ( .B1(n30439), .B2(gray_scale_1[2]), .A1(n15952), .O(n30435)
         );
  OAI12HS U21766 ( .B1(n30446), .B2(gray_scale_1[6]), .A1(n15975), .O(n19935)
         );
  INV1S U21767 ( .I(action_doing[2]), .O(n30413) );
  INV1S U21768 ( .I(medfilt_cnt2_d1[3]), .O(n16050) );
  INV1S U21769 ( .I(medfilt_cnt2_d1[2]), .O(n16051) );
  NR2 U21770 ( .I1(n18537), .I2(n18571), .O(n25372) );
  INV1S U21771 ( .I(cs[0]), .O(n16089) );
  INV1S U21772 ( .I(cs[1]), .O(n18145) );
  INV1S U21773 ( .I(action_doing[0]), .O(n30409) );
  INV1S U21774 ( .I(action_doing[1]), .O(n30410) );
  NR2 U21775 ( .I1(action_doing[0]), .I2(n18458), .O(n19127) );
  AN2B1S U21776 ( .I1(cs_d1[0]), .B1(cs_d1[2]), .O(n30290) );
  AOI22S U21777 ( .A1(medfilt_state_d1[3]), .A2(n16008), .B1(n30290), .B2(
        cs_d1[1]), .O(n16009) );
  NR2 U21778 ( .I1(medfilt_cnt_d1[3]), .I2(n18476), .O(n16049) );
  INV1S U21779 ( .I(medfilt_cnt_d1[0]), .O(n18477) );
  INV1S U21780 ( .I(medfilt_cnt_d1[1]), .O(n18137) );
  NR2 U21781 ( .I1(n18883), .I2(n25050), .O(n25194) );
  INV1S U21782 ( .I(cnt_bdyn_d1[3]), .O(n16053) );
  INV1S U21783 ( .I(cnt_bdyn_d1[2]), .O(n16054) );
  NR2 U21784 ( .I1(n18538), .I2(n18572), .O(n25370) );
  INV1S U21785 ( .I(n30384), .O(n30383) );
  INV1S U21786 ( .I(cnt_dyn_d1[0]), .O(n18478) );
  INV1S U21787 ( .I(cnt_dyn_d1[1]), .O(n18139) );
  AOI22S U21788 ( .A1(n25372), .A2(n25194), .B1(n25370), .B2(n25193), .O(
        n16012) );
  INV1S U21789 ( .I(action_done), .O(n18400) );
  AO13S U21790 ( .B1(n25315), .B2(n18400), .B3(n24901), .A1(n16006), .O(n16011) );
  ND2 U21791 ( .I1(n16012), .I2(n25374), .O(n27222) );
  INV1S U21792 ( .I(gray_img[87]), .O(n16013) );
  INV1S U21793 ( .I(gray_img[215]), .O(n16037) );
  ND2S U21794 ( .I1(n16013), .I2(n16037), .O(n20977) );
  NR2 U21795 ( .I1(gray_img[95]), .I2(gray_img[223]), .O(n20978) );
  INV1S U21796 ( .I(gray_img[95]), .O(n25222) );
  INV1S U21797 ( .I(gray_img[94]), .O(n21141) );
  INV1S U21798 ( .I(gray_img[93]), .O(n16020) );
  INV1S U21799 ( .I(gray_img[92]), .O(n16018) );
  INV1S U21800 ( .I(gray_img[91]), .O(n21534) );
  INV1S U21801 ( .I(gray_img[90]), .O(n16015) );
  FA1S U21802 ( .A(intadd_188_B_0_), .B(intadd_188_A_0_), .CI(gray_img[217]), 
        .CO(n16014) );
  FA1S U21803 ( .A(gray_img[218]), .B(n16015), .CI(n16014), .CO(n16016) );
  FA1S U21804 ( .A(gray_img[219]), .B(n21534), .CI(n16016), .CO(n16017) );
  FA1S U21805 ( .A(gray_img[220]), .B(n16018), .CI(n16017), .CO(n16019) );
  FA1S U21806 ( .A(gray_img[221]), .B(n16020), .CI(n16019), .CO(n16021) );
  NR2 U21807 ( .I1(n25222), .I2(n16022), .O(n16024) );
  AOI12HS U21808 ( .B1(n16022), .B2(n25222), .A1(gray_img[223]), .O(n16023) );
  MXL2HS U21809 ( .A(gray_img[94]), .B(gray_img[222]), .S(n16038), .OB(n26729)
         );
  INV1S U21810 ( .I(gray_img[214]), .O(n16035) );
  INV1S U21811 ( .I(gray_img[213]), .O(n16033) );
  INV1S U21812 ( .I(gray_img[212]), .O(n16031) );
  INV1S U21813 ( .I(gray_img[211]), .O(n16029) );
  INV1S U21814 ( .I(gray_img[210]), .O(n16027) );
  INV1S U21815 ( .I(gray_img[209]), .O(n16025) );
  MXL2HS U21816 ( .A(gray_img[93]), .B(gray_img[221]), .S(n16038), .OB(n26831)
         );
  MXL2HS U21817 ( .A(gray_img[92]), .B(gray_img[220]), .S(n16038), .OB(n16060)
         );
  MXL2HS U21818 ( .A(gray_img[91]), .B(gray_img[219]), .S(n16038), .OB(n16068)
         );
  MUX2S U21819 ( .A(gray_img[210]), .B(gray_img[82]), .S(n23483), .O(n26838)
         );
  MXL2HS U21820 ( .A(gray_img[90]), .B(gray_img[218]), .S(n16038), .OB(n26836)
         );
  MXL2HS U21821 ( .A(gray_img[88]), .B(gray_img[216]), .S(n16038), .OB(n23489)
         );
  MXL2HS U21822 ( .A(gray_img[89]), .B(gray_img[217]), .S(n16038), .OB(n26845)
         );
  MUX2S U21823 ( .A(gray_img[209]), .B(gray_img[81]), .S(n23483), .O(n26848)
         );
  INV1S U21824 ( .I(n16044), .O(n16045) );
  INV1S U21825 ( .I(n26849), .O(n16062) );
  INV1S U21826 ( .I(n16046), .O(n16061) );
  INV1S U21827 ( .I(n27447), .O(n29032) );
  NR2 U21828 ( .I1(n18819), .I2(n25050), .O(n25245) );
  INV1S U21829 ( .I(medfilt_cnt2_d1[0]), .O(n18469) );
  INV1S U21830 ( .I(medfilt_cnt2_d1[1]), .O(n18094) );
  NR2 U21831 ( .I1(n18542), .I2(n18509), .O(n25273) );
  INV1S U21832 ( .I(cnt_bdyn_d1[0]), .O(n18470) );
  INV1S U21833 ( .I(cnt_bdyn_d1[1]), .O(n18095) );
  NR2 U21834 ( .I1(n18543), .I2(n18510), .O(n25271) );
  AOI22S U21835 ( .A1(n25245), .A2(n25273), .B1(n25244), .B2(n25271), .O(
        n16055) );
  MUX2S U21836 ( .A(n29032), .B(n26842), .S(gray_img[44]), .O(n16059) );
  INV1S U21837 ( .I(medfilt_out_reg[4]), .O(n16056) );
  NR2 U21838 ( .I1(n16056), .I2(n18734), .O(n16057) );
  AOI12HS U21839 ( .B1(mem_data_a_out[4]), .B2(n16010), .A1(n16057), .O(n29837) );
  OAI12HS U21840 ( .B1(n16062), .B2(n16061), .A1(n16005), .O(n14244) );
  INV1S U21841 ( .I(n16063), .O(n16069) );
  INV1S U21842 ( .I(medfilt_out_reg[3]), .O(n16064) );
  NR2 U21843 ( .I1(n16064), .I2(n18734), .O(n16065) );
  OAI12HS U21844 ( .B1(n16062), .B2(n16069), .A1(n16004), .O(n14245) );
  INV2 U21845 ( .I(cnt_cro_x[1]), .O(n30375) );
  NR2 U21846 ( .I1(cnt_cro_x[0]), .I2(cnt_cro_3[0]), .O(n16070) );
  OR2P U21847 ( .I1(n30375), .I2(n16070), .O(n16224) );
  ND2S U21848 ( .I1(cnt_cro_x[2]), .I2(cnt_cro_3[1]), .O(n16071) );
  OAI22S U21849 ( .A1(cnt_cro_x[2]), .A2(n16226), .B1(n16224), .B2(n16071), 
        .O(n16235) );
  INV1S U21850 ( .I(cnt_cro_x[3]), .O(n30374) );
  XOR2HS U21851 ( .I1(cnt_dyn_base[2]), .I2(cnt_cro_y[2]), .O(n16073) );
  XOR2HS U21852 ( .I1(cnt_dyn_base[1]), .I2(cnt_cro_y[1]), .O(n16072) );
  NR2 U21853 ( .I1(n16073), .I2(n16072), .O(n16076) );
  XNR2HS U21854 ( .I1(cnt_dyn_base[3]), .I2(cnt_cro_y[3]), .O(n16075) );
  XNR2HS U21855 ( .I1(cnt_dyn_base[0]), .I2(cnt_cro_y[0]), .O(n16074) );
  ND3S U21856 ( .I1(n16076), .I2(n16075), .I3(n16074), .O(n19400) );
  NR2P U21857 ( .I1(cnt_cro_y[1]), .I2(n24948), .O(n16079) );
  OR2P U21858 ( .I1(cnt_cro_3b3[0]), .I2(cnt_cro_y[0]), .O(n16101) );
  INV1 U21859 ( .I(cnt_cro_y[1]), .O(n25038) );
  NR2 U21860 ( .I1(cnt_cro_3b3[1]), .I2(n25038), .O(n16077) );
  NR2P U21861 ( .I1(n16101), .I2(n16077), .O(n16078) );
  NR2F U21862 ( .I1(n16079), .I2(n16078), .O(n16111) );
  INV1S U21863 ( .I(cnt_cro_y[3]), .O(n25045) );
  XOR2HS U21864 ( .I1(cnt_dyn_base[0]), .I2(cnt_cro_x[0]), .O(n16084) );
  XOR2HS U21865 ( .I1(cnt_dyn_base[3]), .I2(cnt_cro_x[3]), .O(n16083) );
  XNR2HS U21866 ( .I1(cnt_dyn_base[1]), .I2(cnt_cro_x[1]), .O(n16081) );
  XNR2HS U21867 ( .I1(cnt_dyn_base[2]), .I2(cnt_cro_x[2]), .O(n16080) );
  ND2S U21868 ( .I1(n16081), .I2(n16080), .O(n16082) );
  NR3 U21869 ( .I1(n16084), .I2(n16083), .I3(n16082), .O(n19402) );
  INV1S U21870 ( .I(cnt_cro_3[1]), .O(n24940) );
  NR2 U21871 ( .I1(cnt_cro_3[0]), .I2(n24940), .O(n19397) );
  ND2S U21872 ( .I1(n19402), .I2(n19397), .O(n16085) );
  OAI112HS U21873 ( .C1(n19396), .C2(n19400), .A1(n16086), .B1(n16085), .O(
        n16087) );
  AOI13HS U21874 ( .B1(n30375), .B2(n16235), .B3(n30374), .A1(n16087), .O(
        n17949) );
  OA13S U21875 ( .B1(cnt_20[1]), .B2(cnt_20[0]), .B3(cnt_20[2]), .A1(cnt_20[3]), .O(n16088) );
  NR3 U21876 ( .I1(cnt_20[5]), .I2(cnt_20[4]), .I3(n16088), .O(n25040) );
  NR2 U21877 ( .I1(n18145), .I2(n24910), .O(n30411) );
  INV1S U21878 ( .I(n30411), .O(n24897) );
  OR2 U21879 ( .I1(n17949), .I2(n17950), .O(n30220) );
  INV1S U21880 ( .I(cro_mac[11]), .O(n17953) );
  INV1S U21881 ( .I(cnt_cro_3b3[0]), .O(n24951) );
  INV1S U21882 ( .I(cnt_cro_3[0]), .O(n16090) );
  NR2 U21883 ( .I1(cnt_cro_3b3[1]), .I2(n24943), .O(n17581) );
  NR2 U21884 ( .I1(cnt_cro_3b3[1]), .I2(n24939), .O(n17579) );
  ND2S U21885 ( .I1(n16091), .I2(cnt_cro_3b3[0]), .O(n16094) );
  NR2 U21886 ( .I1(n24948), .I2(n24940), .O(n17584) );
  NR2 U21887 ( .I1(n24948), .I2(n24943), .O(n17583) );
  AOI22S U21888 ( .A1(n17584), .A2(template_reg[66]), .B1(n17583), .B2(
        template_reg[58]), .O(n16093) );
  NR2 U21889 ( .I1(n24948), .I2(n24939), .O(n17585) );
  ND2S U21890 ( .I1(n17585), .I2(template_reg[50]), .O(n16092) );
  ND2 U21891 ( .I1(n16113), .I2(cnt_cro_y[2]), .O(n16099) );
  XNR2HS U21892 ( .I1(cnt_cro_3b3[1]), .I2(cnt_cro_y[2]), .O(n16097) );
  ND2S U21893 ( .I1(n16111), .I2(n16097), .O(n16098) );
  OAI112HP U21894 ( .C1(n16111), .C2(n16100), .A1(n16099), .B1(n16098), .O(
        n16159) );
  XOR2HS U21895 ( .I1(cnt_cro_3b3[1]), .I2(cnt_cro_y[1]), .O(n16102) );
  NR2 U21896 ( .I1(n16157), .I2(n16154), .O(n16124) );
  ND2P U21897 ( .I1(n16159), .I2(n16124), .O(n16205) );
  OR2 U21898 ( .I1(cnt_cro_3[1]), .I2(n16224), .O(n16105) );
  ND3 U21899 ( .I1(n16103), .I2(n16224), .I3(cnt_cro_3[1]), .O(n16104) );
  ND3P U21900 ( .I1(n16226), .I2(n16105), .I3(n16104), .O(n16231) );
  XOR2HS U21901 ( .I1(cnt_cro_x[0]), .I2(cnt_cro_3[0]), .O(n16106) );
  OAI12HS U21902 ( .B1(n16106), .B2(cnt_dyn_base[0]), .A1(cnt_dyn_base[1]), 
        .O(n16230) );
  INV1S U21903 ( .I(n16106), .O(n16109) );
  NR2P U21904 ( .I1(cnt_dyn_base[0]), .I2(cnt_dyn_base[1]), .O(n18385) );
  ND2 U21905 ( .I1(n16109), .I2(n18385), .O(n16228) );
  ND2S U21906 ( .I1(n16230), .I2(n16228), .O(n16107) );
  ND2 U21907 ( .I1(n16107), .I2(action_5_flag), .O(n16108) );
  XOR2H U21908 ( .I1(n16231), .I2(n16108), .O(n16147) );
  INV1S U21909 ( .I(action_5_flag), .O(n16241) );
  INV2 U21910 ( .I(cnt_dyn_base[0]), .O(n24898) );
  NR2 U21911 ( .I1(n16241), .I2(n24898), .O(n16110) );
  INV1S U21912 ( .I(n16148), .O(n16118) );
  XNR2HS U21913 ( .I1(cnt_cro_y[2]), .I2(cnt_cro_y[3]), .O(n16115) );
  AOI12HS U21914 ( .B1(n16111), .B2(cnt_cro_3b3[1]), .A1(n25037), .O(n16112)
         );
  XNR2H U21915 ( .I1(n16115), .I2(n16114), .O(n16149) );
  ND2P U21916 ( .I1(n16118), .I2(n16149), .O(n16136) );
  INV2 U21917 ( .I(n16154), .O(n16158) );
  NR2 U21918 ( .I1(n16157), .I2(n16158), .O(n16155) );
  INV1S U21919 ( .I(n16155), .O(n16117) );
  OR2P U21920 ( .I1(n16117), .I2(n16159), .O(n16198) );
  INV2 U21921 ( .I(n16149), .O(n16152) );
  ND2 U21922 ( .I1(n16152), .I2(n16118), .O(n16128) );
  OR2T U21923 ( .I1(n16147), .I2(n16128), .O(n16196) );
  AOI22S U21924 ( .A1(n16116), .A2(gray_img[511]), .B1(n15914), .B2(
        gray_img[1791]), .O(n16133) );
  INV1S U21925 ( .I(n16157), .O(n16120) );
  ND2P U21926 ( .I1(n16126), .I2(n16154), .O(n16164) );
  NR2 U21927 ( .I1(n16164), .I2(n16209), .O(n16121) );
  INV2 U21928 ( .I(n16164), .O(n16140) );
  ND3HT U21929 ( .I1(n16152), .I2(n16135), .I3(n16148), .O(n16207) );
  AOI22S U21930 ( .A1(n17703), .A2(gray_img[639]), .B1(n17767), .B2(
        gray_img[1655]), .O(n16132) );
  ND3HT U21931 ( .I1(n16149), .I2(n16135), .I3(n16148), .O(n16213) );
  NR2 U21932 ( .I1(n16213), .I2(n16205), .O(n16123) );
  INV2 U21933 ( .I(n16123), .O(n17221) );
  INV1S U21934 ( .I(n17221), .O(n16345) );
  INV1S U21935 ( .I(n16124), .O(n16125) );
  NR2 U21936 ( .I1(n16210), .I2(n16196), .O(n16301) );
  AOI22S U21937 ( .A1(n16345), .A2(gray_img[503]), .B1(n15873), .B2(
        gray_img[2047]), .O(n16131) );
  INV2 U21938 ( .I(n15917), .O(n17766) );
  INV1S U21939 ( .I(gray_img[887]), .O(n26387) );
  OR2T U21940 ( .I1(n16135), .I2(n16128), .O(n16204) );
  NR2 U21941 ( .I1(n16168), .I2(n16204), .O(n16129) );
  MOAI1S U21942 ( .A1(n17766), .A2(n26387), .B1(n17765), .B2(gray_img[1903]), 
        .O(n16130) );
  AN4B1S U21943 ( .I1(n16133), .I2(n16132), .I3(n16131), .B1(n16130), .O(
        n16181) );
  AOI22S U21944 ( .A1(n15898), .A2(gray_img[895]), .B1(n15911), .B2(
        gray_img[1919]), .O(n16146) );
  INV1S U21945 ( .I(n16213), .O(n16138) );
  AOI22S U21946 ( .A1(n16137), .A2(gray_img[879]), .B1(n17744), .B2(
        gray_img[631]), .O(n16145) );
  NR2 U21947 ( .I1(n16164), .I2(n16203), .O(n16139) );
  AOI22S U21948 ( .A1(n15948), .A2(gray_img[1911]), .B1(n17709), .B2(
        gray_img[623]), .O(n16144) );
  INV1S U21949 ( .I(n16204), .O(n16141) );
  INV1S U21950 ( .I(gray_img[1647]), .O(n25792) );
  MOAI1S U21951 ( .A1(n17381), .A2(n25792), .B1(n15908), .B2(gray_img[1663]), 
        .O(n16143) );
  OR2P U21952 ( .I1(n16149), .I2(n16151), .O(n16173) );
  NR2 U21953 ( .I1(n16205), .I2(n16174), .O(n16153) );
  AOI22S U21954 ( .A1(n15913), .A2(gray_img[1511]), .B1(n17750), .B2(
        gray_img[487]), .O(n16163) );
  ND3P U21955 ( .I1(n16159), .I2(n16157), .I3(n16154), .O(n16208) );
  AOI22S U21956 ( .A1(n16000), .A2(gray_img[1127]), .B1(n17751), .B2(
        gray_img[1639]), .O(n16162) );
  ND2P U21957 ( .I1(n16159), .I2(n16155), .O(n16212) );
  ND3P U21958 ( .I1(n16159), .I2(n16158), .I3(n16157), .O(n16211) );
  AOI22S U21959 ( .A1(n15909), .A2(gray_img[231]), .B1(gray_img[1383]), .B2(
        n15903), .O(n16161) );
  OR2P U21960 ( .I1(n16210), .I2(n16173), .O(n17753) );
  INV1S U21961 ( .I(gray_img[2023]), .O(n25848) );
  MOAI1S U21962 ( .A1(n17753), .A2(n25848), .B1(n17752), .B2(gray_img[359]), 
        .O(n16160) );
  AN4B1S U21963 ( .I1(n16163), .I2(n16162), .I3(n16161), .B1(n16160), .O(
        n16179) );
  NR2T U21964 ( .I1(n16164), .I2(n16174), .O(n16165) );
  INV1S U21965 ( .I(gray_img[615]), .O(n26174) );
  NR2 U21966 ( .I1(n16168), .I2(n16174), .O(n16166) );
  NR2 U21967 ( .I1(n16212), .I2(n16173), .O(n16167) );
  INV2 U21968 ( .I(n17759), .O(n17518) );
  INV1S U21969 ( .I(gray_img[1255]), .O(n28043) );
  MOAI1S U21970 ( .A1(n17518), .A2(n28043), .B1(n15901), .B2(gray_img[1895]), 
        .O(n16169) );
  NR2 U21971 ( .I1(n16170), .I2(n16169), .O(n16177) );
  INV1S U21972 ( .I(n16174), .O(n16172) );
  INV1S U21973 ( .I(n16198), .O(n16171) );
  INV3 U21974 ( .I(n17760), .O(n17639) );
  AOI22S U21975 ( .A1(n15900), .A2(gray_img[999]), .B1(n17639), .B2(
        gray_img[743]), .O(n16176) );
  INV2 U21976 ( .I(n16461), .O(n17478) );
  AOI22S U21977 ( .A1(n15902), .A2(gray_img[1767]), .B1(n17478), .B2(
        gray_img[103]), .O(n16175) );
  ND3S U21978 ( .I1(n16177), .I2(n16176), .I3(n16175), .O(n16178) );
  AN4B1S U21979 ( .I1(n16181), .I2(n16180), .I3(n16179), .B1(n16178), .O(
        n16222) );
  NR2 U21980 ( .I1(n16212), .I2(n16204), .O(n16182) );
  AOI22S U21981 ( .A1(n15872), .A2(gray_img[1151]), .B1(n17785), .B2(
        gray_img[1263]), .O(n16187) );
  NR2 U21982 ( .I1(n16212), .I2(n16203), .O(n16183) );
  AOI22S U21983 ( .A1(n15878), .A2(gray_img[1399]), .B1(n17787), .B2(
        gray_img[239]), .O(n16186) );
  AOI22S U21984 ( .A1(n17137), .A2(gray_img[119]), .B1(n15949), .B2(
        gray_img[1527]), .O(n16185) );
  INV1S U21985 ( .I(gray_img[2031]), .O(n25860) );
  MOAI1S U21986 ( .A1(n15894), .A2(n25860), .B1(n17786), .B2(gray_img[767]), 
        .O(n16184) );
  AN4B1S U21987 ( .I1(n16187), .I2(n16186), .I3(n16185), .B1(n16184), .O(
        n16195) );
  AOI22S U21988 ( .A1(n15876), .A2(gray_img[1783]), .B1(n16188), .B2(
        gray_img[1279]), .O(n16194) );
  NR2 U21989 ( .I1(n16205), .I2(n16203), .O(n16189) );
  AOI22S U21990 ( .A1(n17778), .A2(gray_img[495]), .B1(n15895), .B2(
        gray_img[1535]), .O(n16193) );
  NR2 U21991 ( .I1(n16211), .I2(n16209), .O(n17197) );
  AOI22S U21992 ( .A1(n17780), .A2(gray_img[383]), .B1(gray_img[111]), .B2(
        n17779), .O(n16191) );
  NR2P U21993 ( .I1(n16198), .I2(n16203), .O(n16368) );
  AOI22S U21994 ( .A1(n15877), .A2(gray_img[367]), .B1(n15899), .B2(
        gray_img[751]), .O(n16190) );
  ND2S U21995 ( .I1(n16191), .I2(n16190), .O(n16192) );
  AN4B1S U21996 ( .I1(n16195), .I2(n16194), .I3(n16193), .B1(n16192), .O(
        n16221) );
  NR2 U21997 ( .I1(n16211), .I2(n16196), .O(n16197) );
  BUF2 U21998 ( .I(n16197), .O(n16531) );
  INV2 U21999 ( .I(n16531), .O(n16668) );
  AOI22S U22000 ( .A1(n15874), .A2(gray_img[1135]), .B1(n16531), .B2(
        gray_img[1407]), .O(n16202) );
  AOI22S U22001 ( .A1(n16001), .A2(gray_img[759]), .B1(n15875), .B2(
        gray_img[127]), .O(n16201) );
  NR2 U22002 ( .I1(n16210), .I2(n16213), .O(n16380) );
  AOI22S U22003 ( .A1(n17807), .A2(gray_img[1015]), .B1(n15951), .B2(
        gray_img[1271]), .O(n16200) );
  NR2 U22004 ( .I1(n16212), .I2(n16209), .O(n16280) );
  INV1S U22005 ( .I(gray_img[255]), .O(n27568) );
  MOAI1S U22006 ( .A1(n17533), .A2(n27568), .B1(n17805), .B2(gray_img[1775]), 
        .O(n16199) );
  AN4B1S U22007 ( .I1(n16202), .I2(n16201), .I3(n16200), .B1(n16199), .O(
        n16219) );
  OR2P U22008 ( .I1(n16210), .I2(n16203), .O(n17718) );
  INV1 U22009 ( .I(n17718), .O(n17795) );
  AOI22S U22010 ( .A1(n17796), .A2(gray_img[1391]), .B1(n17795), .B2(
        gray_img[1007]), .O(n16218) );
  NR2P U22011 ( .I1(n16210), .I2(n16207), .O(n17716) );
  NR2 U22012 ( .I1(n16205), .I2(n16204), .O(n16206) );
  AOI22S U22013 ( .A1(n15897), .A2(gray_img[2039]), .B1(n17797), .B2(
        gray_img[1519]), .O(n16217) );
  NR2 U22014 ( .I1(n16210), .I2(n16209), .O(n16325) );
  AOI22S U22015 ( .A1(n17605), .A2(gray_img[1143]), .B1(n15879), .B2(
        gray_img[1023]), .O(n16215) );
  NR2P U22016 ( .I1(n16211), .I2(n16213), .O(n17798) );
  AOI22S U22017 ( .A1(n17798), .A2(gray_img[375]), .B1(n15950), .B2(
        gray_img[247]), .O(n16214) );
  ND2S U22018 ( .I1(n16215), .I2(n16214), .O(n16216) );
  AN4B1S U22019 ( .I1(n16219), .I2(n16218), .I3(n16217), .B1(n16216), .O(
        n16220) );
  NR2 U22020 ( .I1(n24940), .I2(n16224), .O(n16223) );
  NR2 U22021 ( .I1(cnt_cro_x[2]), .I2(n16223), .O(n16227) );
  OAI12HS U22022 ( .B1(n24940), .B2(n16224), .A1(n16226), .O(n16225) );
  AOI22S U22023 ( .A1(n16227), .A2(n16226), .B1(n16225), .B2(cnt_cro_x[2]), 
        .O(n16237) );
  INV1S U22024 ( .I(n16237), .O(n16234) );
  INV1S U22025 ( .I(n16228), .O(n16229) );
  AOI12HS U22026 ( .B1(n16231), .B2(n16230), .A1(n16229), .O(n16236) );
  XOR2HS U22027 ( .I1(cnt_dyn_base[2]), .I2(n16236), .O(n16232) );
  NR2 U22028 ( .I1(n16241), .I2(n16232), .O(n16233) );
  XNR2HS U22029 ( .I1(n16234), .I2(n16233), .O(n16340) );
  INV1S U22030 ( .I(n16340), .O(n16391) );
  XOR2HS U22031 ( .I1(cnt_cro_x[3]), .I2(n16235), .O(n16243) );
  NR2 U22032 ( .I1(cnt_dyn_base[2]), .I2(n16236), .O(n16238) );
  MOAI1S U22033 ( .A1(n16238), .A2(n16237), .B1(cnt_dyn_base[2]), .B2(n16236), 
        .O(n16239) );
  XOR2HS U22034 ( .I1(cnt_dyn_base[3]), .I2(n16239), .O(n16240) );
  NR2 U22035 ( .I1(n16241), .I2(n16240), .O(n16242) );
  XNR2HS U22036 ( .I1(n16243), .I2(n16242), .O(n16339) );
  INV4 U22037 ( .I(n17381), .O(n17743) );
  AOI22S U22038 ( .A1(gray_img[1567]), .A2(n15908), .B1(n17743), .B2(
        gray_img[1551]), .O(n16247) );
  AOI22S U22039 ( .A1(n15898), .A2(gray_img[799]), .B1(n15911), .B2(
        gray_img[1823]), .O(n16246) );
  AOI22S U22040 ( .A1(n15948), .A2(gray_img[1815]), .B1(n17709), .B2(
        gray_img[527]), .O(n16245) );
  INV1S U22041 ( .I(gray_img[535]), .O(n29062) );
  MOAI1S U22042 ( .A1(n17505), .A2(n29062), .B1(n16137), .B2(gray_img[783]), 
        .O(n16244) );
  AN4B1S U22043 ( .I1(n16247), .I2(n16246), .I3(n16245), .B1(n16244), .O(
        n16264) );
  AOI22S U22044 ( .A1(n16116), .A2(gray_img[415]), .B1(gray_img[1695]), .B2(
        n15914), .O(n16251) );
  AOI22S U22045 ( .A1(n17703), .A2(gray_img[543]), .B1(n17767), .B2(
        gray_img[1559]), .O(n16250) );
  AOI22S U22046 ( .A1(n15917), .A2(gray_img[791]), .B1(n17765), .B2(
        gray_img[1807]), .O(n16249) );
  INV1S U22047 ( .I(gray_img[407]), .O(n28746) );
  MOAI1S U22048 ( .A1(n17221), .A2(n28746), .B1(n15873), .B2(gray_img[1951]), 
        .O(n16248) );
  AN4B1S U22049 ( .I1(n16251), .I2(n16250), .I3(n16249), .B1(n16248), .O(
        n16263) );
  INV2 U22050 ( .I(n17753), .O(n17696) );
  AOI22S U22051 ( .A1(n17752), .A2(gray_img[263]), .B1(n17696), .B2(
        gray_img[1927]), .O(n16255) );
  AOI22S U22052 ( .A1(n15913), .A2(gray_img[1415]), .B1(n17750), .B2(
        gray_img[391]), .O(n16254) );
  AOI22S U22053 ( .A1(n15909), .A2(gray_img[135]), .B1(n15903), .B2(
        gray_img[1287]), .O(n16253) );
  INV1S U22054 ( .I(gray_img[1543]), .O(n26600) );
  MOAI1S U22055 ( .A1(n15942), .A2(n26600), .B1(n16000), .B2(gray_img[1031]), 
        .O(n16252) );
  AN4B1S U22056 ( .I1(n16255), .I2(n16254), .I3(n16253), .B1(n16252), .O(
        n16262) );
  INV1S U22057 ( .I(gray_img[519]), .O(n29929) );
  MOAI1S U22058 ( .A1(n17640), .A2(n29929), .B1(n17758), .B2(gray_img[775]), 
        .O(n16257) );
  INV1S U22059 ( .I(gray_img[1159]), .O(n26639) );
  MOAI1S U22060 ( .A1(n17518), .A2(n26639), .B1(n15901), .B2(gray_img[1799]), 
        .O(n16256) );
  NR2 U22061 ( .I1(n16257), .I2(n16256), .O(n16260) );
  AOI22S U22062 ( .A1(n15900), .A2(gray_img[903]), .B1(n17639), .B2(
        gray_img[647]), .O(n16259) );
  AOI22S U22063 ( .A1(n15902), .A2(gray_img[1671]), .B1(n15912), .B2(
        gray_img[7]), .O(n16258) );
  ND3S U22064 ( .I1(n16260), .I2(n16259), .I3(n16258), .O(n16261) );
  AN4B1S U22065 ( .I1(n16264), .I2(n16263), .I3(n16262), .B1(n16261), .O(
        n16289) );
  AOI22S U22066 ( .A1(n17778), .A2(gray_img[399]), .B1(n15895), .B2(
        gray_img[1439]), .O(n16269) );
  AOI22S U22067 ( .A1(n17591), .A2(gray_img[287]), .B1(n17779), .B2(
        gray_img[15]), .O(n16268) );
  AOI22S U22068 ( .A1(n15876), .A2(gray_img[1687]), .B1(n16188), .B2(
        gray_img[1183]), .O(n16267) );
  INV1S U22069 ( .I(gray_img[271]), .O(n21799) );
  MOAI1S U22070 ( .A1(n16518), .A2(n21799), .B1(n15899), .B2(gray_img[655]), 
        .O(n16266) );
  AN4B1S U22071 ( .I1(n16269), .I2(n16268), .I3(n16267), .B1(n16266), .O(
        n16275) );
  AOI22S U22072 ( .A1(n15872), .A2(gray_img[1055]), .B1(n17785), .B2(
        gray_img[1167]), .O(n16274) );
  AOI22S U22073 ( .A1(gray_img[671]), .A2(n17786), .B1(n15866), .B2(
        gray_img[1935]), .O(n16273) );
  AOI22S U22074 ( .A1(n15878), .A2(gray_img[1303]), .B1(n17787), .B2(
        gray_img[143]), .O(n16271) );
  AOI22S U22075 ( .A1(n17137), .A2(gray_img[23]), .B1(n15949), .B2(
        gray_img[1431]), .O(n16270) );
  ND2S U22076 ( .I1(n16271), .I2(n16270), .O(n16272) );
  AN4B1S U22077 ( .I1(n16275), .I2(n16274), .I3(n16273), .B1(n16272), .O(
        n16288) );
  AOI22S U22078 ( .A1(n17716), .A2(gray_img[1943]), .B1(n17797), .B2(
        gray_img[1423]), .O(n16279) );
  AOI22S U22079 ( .A1(n17605), .A2(gray_img[1047]), .B1(n15879), .B2(
        gray_img[927]), .O(n16278) );
  AOI22S U22080 ( .A1(n17717), .A2(gray_img[279]), .B1(n15950), .B2(
        gray_img[151]), .O(n16277) );
  INV1S U22081 ( .I(gray_img[911]), .O(n29616) );
  MOAI1S U22082 ( .A1(n17718), .A2(n29616), .B1(n17796), .B2(gray_img[1295]), 
        .O(n16276) );
  AN4B1S U22083 ( .I1(n16279), .I2(n16278), .I3(n16277), .B1(n16276), .O(
        n16286) );
  AOI22S U22084 ( .A1(n16001), .A2(gray_img[663]), .B1(n15896), .B2(
        gray_img[31]), .O(n16285) );
  AOI22S U22085 ( .A1(n17723), .A2(gray_img[1039]), .B1(n16531), .B2(
        gray_img[1311]), .O(n16284) );
  AOI22S U22086 ( .A1(n17806), .A2(gray_img[159]), .B1(n17805), .B2(
        gray_img[1679]), .O(n16282) );
  AOI22S U22087 ( .A1(n17807), .A2(gray_img[919]), .B1(n15951), .B2(
        gray_img[1175]), .O(n16281) );
  ND2S U22088 ( .I1(n16282), .I2(n16281), .O(n16283) );
  AN4B1S U22089 ( .I1(n16286), .I2(n16285), .I3(n16284), .B1(n16283), .O(
        n16287) );
  ND3S U22090 ( .I1(n16289), .I2(n16288), .I3(n16287), .O(n16290) );
  INV1S U22091 ( .I(n16339), .O(n16390) );
  AOI22S U22092 ( .A1(n16291), .A2(n17819), .B1(n16290), .B2(n17688), .O(
        n16395) );
  AOI22S U22093 ( .A1(n15913), .A2(gray_img[1479]), .B1(n17750), .B2(
        gray_img[455]), .O(n16295) );
  AOI22S U22094 ( .A1(n16000), .A2(gray_img[1095]), .B1(n17751), .B2(
        gray_img[1607]), .O(n16294) );
  AOI22S U22095 ( .A1(n15909), .A2(gray_img[199]), .B1(gray_img[1351]), .B2(
        n15903), .O(n16293) );
  INV1S U22096 ( .I(gray_img[1991]), .O(n23560) );
  MOAI1S U22097 ( .A1(n17753), .A2(n23560), .B1(n17752), .B2(gray_img[327]), 
        .O(n16292) );
  AN4B1S U22098 ( .I1(n16295), .I2(n16294), .I3(n16293), .B1(n16292), .O(
        n16314) );
  AOI22S U22099 ( .A1(n15902), .A2(gray_img[1735]), .B1(n17478), .B2(
        gray_img[71]), .O(n16300) );
  AOI22S U22100 ( .A1(n17758), .A2(gray_img[839]), .B1(n16165), .B2(
        gray_img[583]), .O(n16299) );
  AOI22S U22101 ( .A1(n17759), .A2(gray_img[1223]), .B1(n15901), .B2(
        gray_img[1863]), .O(n16298) );
  INV1S U22102 ( .I(gray_img[711]), .O(n27146) );
  MOAI1S U22103 ( .A1(n17760), .A2(n27146), .B1(n15900), .B2(gray_img[967]), 
        .O(n16297) );
  AN4B1S U22104 ( .I1(n16300), .I2(n16299), .I3(n16298), .B1(n16297), .O(
        n16313) );
  AOI22S U22105 ( .A1(n16116), .A2(gray_img[479]), .B1(n15914), .B2(
        gray_img[1759]), .O(n16305) );
  AOI22S U22106 ( .A1(n16345), .A2(gray_img[471]), .B1(n15873), .B2(
        gray_img[2015]), .O(n16304) );
  AOI22S U22107 ( .A1(n15917), .A2(gray_img[855]), .B1(n17765), .B2(
        gray_img[1871]), .O(n16303) );
  INV1S U22108 ( .I(gray_img[1623]), .O(n25524) );
  MOAI1S U22109 ( .A1(n17704), .A2(n25524), .B1(n17703), .B2(gray_img[607]), 
        .O(n16302) );
  AN4B1S U22110 ( .I1(n16305), .I2(n16304), .I3(n16303), .B1(n16302), .O(
        n16312) );
  INV1S U22111 ( .I(gray_img[599]), .O(n27025) );
  MOAI1S U22112 ( .A1(n17505), .A2(n27025), .B1(n16137), .B2(gray_img[847]), 
        .O(n16307) );
  INV1S U22113 ( .I(gray_img[1615]), .O(n25666) );
  MOAI1S U22114 ( .A1(n17381), .A2(n25666), .B1(n15908), .B2(gray_img[1631]), 
        .O(n16306) );
  NR2 U22115 ( .I1(n16307), .I2(n16306), .O(n16310) );
  AOI22S U22116 ( .A1(n15898), .A2(gray_img[863]), .B1(n15911), .B2(
        gray_img[1887]), .O(n16309) );
  AOI22S U22117 ( .A1(n15948), .A2(gray_img[1879]), .B1(n17709), .B2(
        gray_img[591]), .O(n16308) );
  ND3S U22118 ( .I1(n16310), .I2(n16309), .I3(n16308), .O(n16311) );
  AN4B1S U22119 ( .I1(n16314), .I2(n16313), .I3(n16312), .B1(n16311), .O(
        n16338) );
  AOI22S U22120 ( .A1(n15872), .A2(gray_img[1119]), .B1(n17785), .B2(
        gray_img[1231]), .O(n16318) );
  AOI22S U22121 ( .A1(n15878), .A2(gray_img[1367]), .B1(n17787), .B2(
        gray_img[207]), .O(n16317) );
  AOI22S U22122 ( .A1(n17137), .A2(gray_img[87]), .B1(n15949), .B2(
        gray_img[1495]), .O(n16316) );
  INV1S U22123 ( .I(gray_img[1999]), .O(n25001) );
  MOAI1S U22124 ( .A1(n15894), .A2(n25001), .B1(n17786), .B2(gray_img[735]), 
        .O(n16315) );
  AN4B1S U22125 ( .I1(n16318), .I2(n16317), .I3(n16316), .B1(n16315), .O(
        n16324) );
  AOI22S U22126 ( .A1(n15876), .A2(gray_img[1751]), .B1(n16188), .B2(
        gray_img[1247]), .O(n16323) );
  AOI22S U22127 ( .A1(n17778), .A2(gray_img[463]), .B1(n15895), .B2(
        gray_img[1503]), .O(n16322) );
  AOI22S U22128 ( .A1(n17591), .A2(gray_img[351]), .B1(n17779), .B2(
        gray_img[79]), .O(n16320) );
  AOI22S U22129 ( .A1(n15877), .A2(gray_img[335]), .B1(n15899), .B2(
        gray_img[719]), .O(n16319) );
  ND2S U22130 ( .I1(n16320), .I2(n16319), .O(n16321) );
  AN4B1S U22131 ( .I1(n16324), .I2(n16323), .I3(n16322), .B1(n16321), .O(
        n16337) );
  AOI22S U22132 ( .A1(gray_img[2007]), .A2(n15897), .B1(n17797), .B2(
        gray_img[1487]), .O(n16329) );
  AOI22S U22133 ( .A1(n17605), .A2(gray_img[1111]), .B1(n15879), .B2(
        gray_img[991]), .O(n16328) );
  AOI22S U22134 ( .A1(n17717), .A2(gray_img[343]), .B1(n15950), .B2(
        gray_img[215]), .O(n16327) );
  INV1S U22135 ( .I(gray_img[975]), .O(n22982) );
  MOAI1S U22136 ( .A1(n17718), .A2(n22982), .B1(n17796), .B2(gray_img[1359]), 
        .O(n16326) );
  AN4B1S U22137 ( .I1(n16329), .I2(n16328), .I3(n16327), .B1(n16326), .O(
        n16335) );
  AOI22S U22138 ( .A1(n16001), .A2(gray_img[727]), .B1(n15875), .B2(
        gray_img[95]), .O(n16334) );
  INV1 U22139 ( .I(n16379), .O(n17723) );
  AOI22S U22140 ( .A1(n17723), .A2(gray_img[1103]), .B1(n16531), .B2(
        gray_img[1375]), .O(n16333) );
  AOI22S U22141 ( .A1(n17806), .A2(gray_img[223]), .B1(n17805), .B2(
        gray_img[1743]), .O(n16331) );
  AOI22S U22142 ( .A1(n17807), .A2(gray_img[983]), .B1(n15951), .B2(
        gray_img[1239]), .O(n16330) );
  ND2S U22143 ( .I1(n16331), .I2(n16330), .O(n16332) );
  AN4B1S U22144 ( .I1(n16335), .I2(n16334), .I3(n16333), .B1(n16332), .O(
        n16336) );
  ND3S U22145 ( .I1(n16338), .I2(n16337), .I3(n16336), .O(n16393) );
  AOI22S U22146 ( .A1(n15908), .A2(gray_img[1599]), .B1(n17743), .B2(
        gray_img[1583]), .O(n16344) );
  AOI22S U22147 ( .A1(n15898), .A2(gray_img[831]), .B1(n15911), .B2(
        gray_img[1855]), .O(n16343) );
  AOI22S U22148 ( .A1(n16137), .A2(gray_img[815]), .B1(n17744), .B2(
        gray_img[567]), .O(n16342) );
  INV1S U22149 ( .I(gray_img[559]), .O(n28619) );
  MOAI1S U22150 ( .A1(n17745), .A2(n28619), .B1(n15948), .B2(gray_img[1847]), 
        .O(n16341) );
  AN4B1S U22151 ( .I1(n16344), .I2(n16343), .I3(n16342), .B1(n16341), .O(
        n16362) );
  AOI22S U22152 ( .A1(n16116), .A2(gray_img[447]), .B1(n15914), .B2(
        gray_img[1727]), .O(n16349) );
  AOI22S U22153 ( .A1(n17703), .A2(gray_img[575]), .B1(n17767), .B2(
        gray_img[1591]), .O(n16348) );
  AOI22S U22154 ( .A1(n16345), .A2(gray_img[439]), .B1(n15873), .B2(
        gray_img[1983]), .O(n16347) );
  INV1S U22155 ( .I(gray_img[823]), .O(n26110) );
  MOAI1S U22156 ( .A1(n17766), .A2(n26110), .B1(n17765), .B2(gray_img[1839]), 
        .O(n16346) );
  AN4B1S U22157 ( .I1(n16349), .I2(n16348), .I3(n16347), .B1(n16346), .O(
        n16361) );
  AOI22S U22158 ( .A1(n15913), .A2(gray_img[1447]), .B1(n17750), .B2(
        gray_img[423]), .O(n16353) );
  AOI22S U22159 ( .A1(n16000), .A2(gray_img[1063]), .B1(n17751), .B2(
        gray_img[1575]), .O(n16352) );
  AOI22S U22160 ( .A1(n15909), .A2(gray_img[167]), .B1(n15903), .B2(
        gray_img[1319]), .O(n16351) );
  INV1S U22161 ( .I(gray_img[1959]), .O(n26668) );
  MOAI1S U22162 ( .A1(n17753), .A2(n26668), .B1(n17752), .B2(gray_img[295]), 
        .O(n16350) );
  AN4B1S U22163 ( .I1(n16353), .I2(n16352), .I3(n16351), .B1(n16350), .O(
        n16360) );
  INV1S U22164 ( .I(gray_img[551]), .O(n28632) );
  MOAI1S U22165 ( .A1(n17640), .A2(n28632), .B1(n17758), .B2(gray_img[807]), 
        .O(n16355) );
  INV1S U22166 ( .I(gray_img[1191]), .O(n23020) );
  MOAI1S U22167 ( .A1(n17518), .A2(n23020), .B1(n15901), .B2(gray_img[1831]), 
        .O(n16354) );
  NR2 U22168 ( .I1(n16355), .I2(n16354), .O(n16358) );
  AOI22S U22169 ( .A1(n15900), .A2(gray_img[935]), .B1(n17639), .B2(
        gray_img[679]), .O(n16357) );
  AOI22S U22170 ( .A1(n15902), .A2(gray_img[1703]), .B1(n15912), .B2(
        gray_img[39]), .O(n16356) );
  ND3S U22171 ( .I1(n16358), .I2(n16357), .I3(n16356), .O(n16359) );
  AN4B1S U22172 ( .I1(n16362), .I2(n16361), .I3(n16360), .B1(n16359), .O(
        n16389) );
  AOI22S U22173 ( .A1(n15872), .A2(gray_img[1087]), .B1(n17785), .B2(
        gray_img[1199]), .O(n16367) );
  AOI22S U22174 ( .A1(gray_img[1335]), .A2(n15878), .B1(n17787), .B2(
        gray_img[175]), .O(n16366) );
  AOI22S U22175 ( .A1(n17137), .A2(gray_img[55]), .B1(n15949), .B2(
        gray_img[1463]), .O(n16365) );
  INV1S U22176 ( .I(gray_img[1967]), .O(n26681) );
  MOAI1S U22177 ( .A1(n15894), .A2(n26681), .B1(n17786), .B2(gray_img[703]), 
        .O(n16364) );
  AN4B1S U22178 ( .I1(n16367), .I2(n16366), .I3(n16365), .B1(n16364), .O(
        n16374) );
  AOI22S U22179 ( .A1(n15876), .A2(gray_img[1719]), .B1(n16188), .B2(
        gray_img[1215]), .O(n16373) );
  AOI22S U22180 ( .A1(n17778), .A2(gray_img[431]), .B1(n15895), .B2(
        gray_img[1471]), .O(n16372) );
  AOI22S U22181 ( .A1(n17780), .A2(gray_img[319]), .B1(n17779), .B2(
        gray_img[47]), .O(n16370) );
  AOI22S U22182 ( .A1(n15877), .A2(gray_img[303]), .B1(n16368), .B2(
        gray_img[687]), .O(n16369) );
  ND2S U22183 ( .I1(n16370), .I2(n16369), .O(n16371) );
  AN4B1S U22184 ( .I1(n16374), .I2(n16373), .I3(n16372), .B1(n16371), .O(
        n16388) );
  AOI22S U22185 ( .A1(n15897), .A2(gray_img[1975]), .B1(n17797), .B2(
        gray_img[1455]), .O(n16378) );
  AOI22S U22186 ( .A1(n17605), .A2(gray_img[1079]), .B1(n15879), .B2(
        gray_img[959]), .O(n16377) );
  AOI22S U22187 ( .A1(n17717), .A2(gray_img[311]), .B1(n15950), .B2(
        gray_img[183]), .O(n16376) );
  INV1S U22188 ( .I(gray_img[943]), .O(n24985) );
  MOAI1S U22189 ( .A1(n17718), .A2(n24985), .B1(n17796), .B2(gray_img[1327]), 
        .O(n16375) );
  AN4B1S U22190 ( .I1(n16378), .I2(n16377), .I3(n16376), .B1(n16375), .O(
        n16386) );
  AOI22S U22191 ( .A1(n16001), .A2(gray_img[695]), .B1(n15875), .B2(
        gray_img[63]), .O(n16385) );
  AOI22S U22192 ( .A1(n17723), .A2(gray_img[1071]), .B1(n16531), .B2(
        gray_img[1343]), .O(n16384) );
  AOI22S U22193 ( .A1(n17806), .A2(gray_img[191]), .B1(n17805), .B2(
        gray_img[1711]), .O(n16382) );
  AOI22S U22194 ( .A1(n17807), .A2(gray_img[951]), .B1(n15951), .B2(
        gray_img[1207]), .O(n16381) );
  ND2S U22195 ( .I1(n16382), .I2(n16381), .O(n16383) );
  AN4B1S U22196 ( .I1(n16386), .I2(n16385), .I3(n16384), .B1(n16383), .O(
        n16387) );
  ND3S U22197 ( .I1(n16389), .I2(n16388), .I3(n16387), .O(n16392) );
  AOI22S U22198 ( .A1(n16393), .A2(n17690), .B1(n16392), .B2(n17817), .O(
        n16394) );
  ND2S U22199 ( .I1(n16395), .I2(n16394), .O(n16396) );
  INV2 U22200 ( .I(n16396), .O(n17973) );
  NR2 U22201 ( .I1(n15992), .I2(n17973), .O(n17365) );
  ND2S U22202 ( .I1(n16397), .I2(cnt_cro_3b3[0]), .O(n16400) );
  AOI22S U22203 ( .A1(n17584), .A2(template_reg[67]), .B1(n17583), .B2(
        template_reg[59]), .O(n16399) );
  ND2S U22204 ( .I1(n17585), .I2(template_reg[51]), .O(n16398) );
  AOI22S U22205 ( .A1(gray_img[1566]), .A2(n15908), .B1(n17743), .B2(
        gray_img[1550]), .O(n16406) );
  AOI22S U22206 ( .A1(n15898), .A2(gray_img[798]), .B1(n15911), .B2(
        gray_img[1822]), .O(n16405) );
  AOI22S U22207 ( .A1(n15948), .A2(gray_img[1814]), .B1(n17709), .B2(
        gray_img[526]), .O(n16404) );
  INV1S U22208 ( .I(gray_img[534]), .O(n29060) );
  MOAI1S U22209 ( .A1(n17505), .A2(n29060), .B1(n16137), .B2(gray_img[782]), 
        .O(n16403) );
  AN4B1S U22210 ( .I1(n16406), .I2(n16405), .I3(n16404), .B1(n16403), .O(
        n16423) );
  AOI22S U22211 ( .A1(n16116), .A2(gray_img[414]), .B1(gray_img[1694]), .B2(
        n15914), .O(n16410) );
  AOI22S U22212 ( .A1(n17079), .A2(gray_img[406]), .B1(n15873), .B2(
        gray_img[1950]), .O(n16409) );
  AOI22S U22213 ( .A1(n15917), .A2(gray_img[790]), .B1(n17765), .B2(
        gray_img[1806]), .O(n16408) );
  INV1S U22214 ( .I(gray_img[542]), .O(n29076) );
  INV1 U22215 ( .I(n17703), .O(n17674) );
  MOAI1S U22216 ( .A1(n29076), .A2(n17674), .B1(n17767), .B2(gray_img[1558]), 
        .O(n16407) );
  AN4B1S U22217 ( .I1(n16410), .I2(n16409), .I3(n16408), .B1(n16407), .O(
        n16422) );
  AOI22S U22218 ( .A1(n17752), .A2(gray_img[262]), .B1(n17696), .B2(
        gray_img[1926]), .O(n16414) );
  AOI22S U22219 ( .A1(n15913), .A2(gray_img[1414]), .B1(n17750), .B2(
        gray_img[390]), .O(n16413) );
  AOI22S U22220 ( .A1(n15909), .A2(gray_img[134]), .B1(n15903), .B2(
        gray_img[1286]), .O(n16412) );
  INV1S U22221 ( .I(gray_img[1542]), .O(n26598) );
  MOAI1S U22222 ( .A1(n15942), .A2(n26598), .B1(n16000), .B2(gray_img[1030]), 
        .O(n16411) );
  AN4B1S U22223 ( .I1(n16414), .I2(n16413), .I3(n16412), .B1(n16411), .O(
        n16421) );
  INV1S U22224 ( .I(gray_img[518]), .O(n29927) );
  MOAI1S U22225 ( .A1(n17640), .A2(n29927), .B1(n17758), .B2(gray_img[774]), 
        .O(n16416) );
  INV1S U22226 ( .I(gray_img[1158]), .O(n26637) );
  MOAI1S U22227 ( .A1(n17518), .A2(n26637), .B1(n15901), .B2(gray_img[1798]), 
        .O(n16415) );
  NR2 U22228 ( .I1(n16416), .I2(n16415), .O(n16419) );
  AOI22S U22229 ( .A1(n15900), .A2(gray_img[902]), .B1(n17639), .B2(
        gray_img[646]), .O(n16418) );
  AOI22S U22230 ( .A1(n15902), .A2(gray_img[1670]), .B1(n17478), .B2(
        gray_img[6]), .O(n16417) );
  ND3S U22231 ( .I1(n16419), .I2(n16418), .I3(n16417), .O(n16420) );
  AN4B1S U22232 ( .I1(n16423), .I2(n16422), .I3(n16421), .B1(n16420), .O(
        n16446) );
  AOI22S U22233 ( .A1(n17778), .A2(gray_img[398]), .B1(n15895), .B2(
        gray_img[1438]), .O(n16427) );
  AOI22S U22234 ( .A1(n17591), .A2(gray_img[286]), .B1(n17779), .B2(
        gray_img[14]), .O(n16426) );
  AOI22S U22235 ( .A1(n15876), .A2(gray_img[1686]), .B1(n16188), .B2(
        gray_img[1182]), .O(n16425) );
  INV1S U22236 ( .I(gray_img[270]), .O(n21225) );
  MOAI1S U22237 ( .A1(n16518), .A2(n21225), .B1(n15899), .B2(gray_img[654]), 
        .O(n16424) );
  AN4B1S U22238 ( .I1(n16427), .I2(n16426), .I3(n16425), .B1(n16424), .O(
        n16444) );
  INV2 U22239 ( .I(n16668), .O(n17148) );
  AOI22S U22240 ( .A1(n15874), .A2(gray_img[1038]), .B1(n17148), .B2(
        gray_img[1310]), .O(n16431) );
  AOI22S U22241 ( .A1(n16001), .A2(gray_img[662]), .B1(n15875), .B2(
        gray_img[30]), .O(n16430) );
  AOI22S U22242 ( .A1(n17807), .A2(gray_img[918]), .B1(n15951), .B2(
        gray_img[1174]), .O(n16429) );
  INV1S U22243 ( .I(gray_img[158]), .O(n27874) );
  MOAI1S U22244 ( .A1(n17533), .A2(n27874), .B1(n17805), .B2(gray_img[1678]), 
        .O(n16428) );
  AN4B1S U22245 ( .I1(n16431), .I2(n16430), .I3(n16429), .B1(n16428), .O(
        n16443) );
  AOI22S U22246 ( .A1(n15897), .A2(gray_img[1942]), .B1(n17797), .B2(
        gray_img[1422]), .O(n16435) );
  AOI22S U22247 ( .A1(n17605), .A2(gray_img[1046]), .B1(n15879), .B2(
        gray_img[926]), .O(n16434) );
  AOI22S U22248 ( .A1(n17606), .A2(gray_img[278]), .B1(n15950), .B2(
        gray_img[150]), .O(n16433) );
  INV1S U22249 ( .I(gray_img[910]), .O(n29614) );
  MOAI1S U22250 ( .A1(n17718), .A2(n29614), .B1(n17796), .B2(gray_img[1294]), 
        .O(n16432) );
  AN4B1S U22251 ( .I1(n16435), .I2(n16434), .I3(n16433), .B1(n16432), .O(
        n16442) );
  INV1S U22252 ( .I(gray_img[22]), .O(n27861) );
  MOAI1S U22253 ( .A1(n15941), .A2(n27861), .B1(n15949), .B2(gray_img[1430]), 
        .O(n16437) );
  INV1S U22254 ( .I(gray_img[1302]), .O(n29757) );
  MOAI1S U22255 ( .A1(n15944), .A2(n29757), .B1(n17787), .B2(gray_img[142]), 
        .O(n16436) );
  NR2 U22256 ( .I1(n16437), .I2(n16436), .O(n16440) );
  AOI22S U22257 ( .A1(n15872), .A2(gray_img[1054]), .B1(n17785), .B2(
        gray_img[1166]), .O(n16439) );
  AOI22S U22258 ( .A1(gray_img[670]), .A2(n17786), .B1(n15866), .B2(
        gray_img[1934]), .O(n16438) );
  ND3S U22259 ( .I1(n16440), .I2(n16439), .I3(n16438), .O(n16441) );
  AN4B1S U22260 ( .I1(n16444), .I2(n16443), .I3(n16442), .B1(n16441), .O(
        n16445) );
  ND2S U22261 ( .I1(n16446), .I2(n16445), .O(n16494) );
  AOI22S U22262 ( .A1(n15908), .A2(gray_img[1598]), .B1(n17743), .B2(
        gray_img[1582]), .O(n16450) );
  AOI22S U22263 ( .A1(n15898), .A2(gray_img[830]), .B1(n15911), .B2(
        gray_img[1854]), .O(n16449) );
  AOI22S U22264 ( .A1(n16137), .A2(gray_img[814]), .B1(n17744), .B2(
        gray_img[566]), .O(n16448) );
  INV1S U22265 ( .I(gray_img[558]), .O(n28617) );
  MOAI1S U22266 ( .A1(n17745), .A2(n28617), .B1(n15948), .B2(gray_img[1846]), 
        .O(n16447) );
  AN4B1S U22267 ( .I1(n16450), .I2(n16449), .I3(n16448), .B1(n16447), .O(
        n16468) );
  AOI22S U22268 ( .A1(n16116), .A2(gray_img[446]), .B1(n15914), .B2(
        gray_img[1726]), .O(n16454) );
  AOI22S U22269 ( .A1(n17079), .A2(gray_img[438]), .B1(n15873), .B2(
        gray_img[1982]), .O(n16453) );
  AOI22S U22270 ( .A1(n15917), .A2(gray_img[822]), .B1(n17765), .B2(
        gray_img[1838]), .O(n16452) );
  INV1S U22271 ( .I(gray_img[574]), .O(n28153) );
  MOAI1S U22272 ( .A1(n17674), .A2(n28153), .B1(n17767), .B2(gray_img[1590]), 
        .O(n16451) );
  AN4B1S U22273 ( .I1(n16454), .I2(n16453), .I3(n16452), .B1(n16451), .O(
        n16467) );
  AOI22S U22274 ( .A1(n15913), .A2(gray_img[1446]), .B1(n17750), .B2(
        gray_img[422]), .O(n16458) );
  AOI22S U22275 ( .A1(n16000), .A2(gray_img[1062]), .B1(n17751), .B2(
        gray_img[1574]), .O(n16457) );
  AOI22S U22276 ( .A1(n15909), .A2(gray_img[166]), .B1(n15903), .B2(
        gray_img[1318]), .O(n16456) );
  INV1S U22277 ( .I(gray_img[1958]), .O(n26666) );
  MOAI1S U22278 ( .A1(n17753), .A2(n26666), .B1(n17752), .B2(gray_img[294]), 
        .O(n16455) );
  AN4B1S U22279 ( .I1(n16458), .I2(n16457), .I3(n16456), .B1(n16455), .O(
        n16466) );
  INV1S U22280 ( .I(gray_img[550]), .O(n28630) );
  MOAI1S U22281 ( .A1(n17640), .A2(n28630), .B1(n17758), .B2(gray_img[806]), 
        .O(n16460) );
  INV1S U22282 ( .I(gray_img[1190]), .O(n23018) );
  MOAI1S U22283 ( .A1(n17518), .A2(n23018), .B1(n15901), .B2(gray_img[1830]), 
        .O(n16459) );
  NR2 U22284 ( .I1(n16460), .I2(n16459), .O(n16464) );
  AOI22S U22285 ( .A1(n15900), .A2(gray_img[934]), .B1(n17639), .B2(
        gray_img[678]), .O(n16463) );
  AOI22S U22286 ( .A1(n15902), .A2(gray_img[1702]), .B1(n17478), .B2(
        gray_img[38]), .O(n16462) );
  ND3S U22287 ( .I1(n16464), .I2(n16463), .I3(n16462), .O(n16465) );
  AN4B1S U22288 ( .I1(n16468), .I2(n16467), .I3(n16466), .B1(n16465), .O(
        n16492) );
  AOI22S U22289 ( .A1(n15874), .A2(gray_img[1070]), .B1(n17148), .B2(
        gray_img[1342]), .O(n16472) );
  AOI22S U22290 ( .A1(n17806), .A2(gray_img[190]), .B1(n17805), .B2(
        gray_img[1710]), .O(n16471) );
  AOI22S U22291 ( .A1(n17807), .A2(gray_img[950]), .B1(n15951), .B2(
        gray_img[1206]), .O(n16470) );
  INV1S U22292 ( .I(gray_img[62]), .O(n27719) );
  MOAI1S U22293 ( .A1(n15868), .A2(n27719), .B1(n16001), .B2(gray_img[694]), 
        .O(n16469) );
  AN4B1S U22294 ( .I1(n16472), .I2(n16471), .I3(n16470), .B1(n16469), .O(
        n16490) );
  AOI22S U22295 ( .A1(n15872), .A2(gray_img[1086]), .B1(n17785), .B2(
        gray_img[1198]), .O(n16476) );
  AOI22S U22296 ( .A1(gray_img[1334]), .A2(n15878), .B1(n17787), .B2(
        gray_img[174]), .O(n16475) );
  AOI22S U22297 ( .A1(n17137), .A2(gray_img[54]), .B1(n15949), .B2(
        gray_img[1462]), .O(n16474) );
  INV1S U22298 ( .I(gray_img[1966]), .O(n26679) );
  MOAI1S U22299 ( .A1(n15894), .A2(n26679), .B1(n17786), .B2(gray_img[702]), 
        .O(n16473) );
  AN4B1S U22300 ( .I1(n16476), .I2(n16475), .I3(n16474), .B1(n16473), .O(
        n16489) );
  AOI22S U22301 ( .A1(n15897), .A2(gray_img[1974]), .B1(n17797), .B2(
        gray_img[1454]), .O(n16481) );
  AOI22S U22302 ( .A1(n17605), .A2(gray_img[1078]), .B1(n15879), .B2(
        gray_img[958]), .O(n16480) );
  AOI22S U22303 ( .A1(n17606), .A2(gray_img[310]), .B1(n15950), .B2(
        gray_img[182]), .O(n16479) );
  INV1S U22304 ( .I(gray_img[942]), .O(n23218) );
  MOAI1S U22305 ( .A1(n17718), .A2(n23218), .B1(n17796), .B2(gray_img[1326]), 
        .O(n16478) );
  AN4B1S U22306 ( .I1(n16481), .I2(n16480), .I3(n16479), .B1(n16478), .O(
        n16488) );
  INV1S U22307 ( .I(gray_img[1718]), .O(n29219) );
  MOAI1S U22308 ( .A1(n15947), .A2(n29219), .B1(n16188), .B2(gray_img[1214]), 
        .O(n16483) );
  INV1S U22309 ( .I(gray_img[1470]), .O(n18064) );
  MOAI1S U22310 ( .A1(n15867), .A2(n18064), .B1(n17778), .B2(gray_img[430]), 
        .O(n16482) );
  NR2 U22311 ( .I1(n16483), .I2(n16482), .O(n16486) );
  AOI22S U22312 ( .A1(n17591), .A2(gray_img[318]), .B1(n17779), .B2(
        gray_img[46]), .O(n16485) );
  AOI22S U22313 ( .A1(n15877), .A2(gray_img[302]), .B1(n15899), .B2(
        gray_img[686]), .O(n16484) );
  ND3S U22314 ( .I1(n16486), .I2(n16485), .I3(n16484), .O(n16487) );
  AN4B1S U22315 ( .I1(n16490), .I2(n16489), .I3(n16488), .B1(n16487), .O(
        n16491) );
  ND2S U22316 ( .I1(n16492), .I2(n16491), .O(n16493) );
  AOI22S U22317 ( .A1(n16494), .A2(n17688), .B1(n17817), .B2(n16493), .O(
        n16590) );
  AOI22S U22318 ( .A1(n15913), .A2(gray_img[1478]), .B1(n17750), .B2(
        gray_img[454]), .O(n16499) );
  AOI22S U22319 ( .A1(n16000), .A2(gray_img[1094]), .B1(n17751), .B2(
        gray_img[1606]), .O(n16498) );
  AOI22S U22320 ( .A1(n15909), .A2(gray_img[198]), .B1(n15903), .B2(
        gray_img[1350]), .O(n16497) );
  INV1S U22321 ( .I(gray_img[1990]), .O(n23558) );
  MOAI1S U22322 ( .A1(n17753), .A2(n23558), .B1(n17752), .B2(gray_img[326]), 
        .O(n16496) );
  AN4B1S U22323 ( .I1(n16499), .I2(n16498), .I3(n16497), .B1(n16496), .O(
        n16517) );
  AOI22S U22324 ( .A1(n15902), .A2(gray_img[1734]), .B1(n15912), .B2(
        gray_img[70]), .O(n16504) );
  AOI22S U22325 ( .A1(n17758), .A2(gray_img[838]), .B1(n16165), .B2(
        gray_img[582]), .O(n16503) );
  AOI22S U22326 ( .A1(n17759), .A2(gray_img[1222]), .B1(n15901), .B2(
        gray_img[1862]), .O(n16502) );
  INV1S U22327 ( .I(gray_img[710]), .O(n27144) );
  MOAI1S U22328 ( .A1(n17760), .A2(n27144), .B1(n15900), .B2(gray_img[966]), 
        .O(n16501) );
  AN4B1S U22329 ( .I1(n16504), .I2(n16503), .I3(n16502), .B1(n16501), .O(
        n16516) );
  AOI22S U22330 ( .A1(n16116), .A2(gray_img[478]), .B1(n15914), .B2(
        gray_img[1758]), .O(n16508) );
  AOI22S U22331 ( .A1(n17079), .A2(gray_img[470]), .B1(n15873), .B2(
        gray_img[2014]), .O(n16507) );
  AOI22S U22332 ( .A1(n15917), .A2(gray_img[854]), .B1(n17765), .B2(
        gray_img[1870]), .O(n16506) );
  INV1S U22333 ( .I(gray_img[1622]), .O(n25522) );
  MOAI1S U22334 ( .A1(n17704), .A2(n25522), .B1(n17703), .B2(gray_img[606]), 
        .O(n16505) );
  AN4B1S U22335 ( .I1(n16508), .I2(n16507), .I3(n16506), .B1(n16505), .O(
        n16515) );
  INV1S U22336 ( .I(gray_img[598]), .O(n27023) );
  MOAI1S U22337 ( .A1(n17505), .A2(n27023), .B1(n16137), .B2(gray_img[846]), 
        .O(n16510) );
  INV1S U22338 ( .I(gray_img[1614]), .O(n25664) );
  MOAI1S U22339 ( .A1(n17381), .A2(n25664), .B1(n15908), .B2(gray_img[1630]), 
        .O(n16509) );
  NR2 U22340 ( .I1(n16510), .I2(n16509), .O(n16513) );
  AOI22S U22341 ( .A1(n15898), .A2(gray_img[862]), .B1(n15911), .B2(
        gray_img[1886]), .O(n16512) );
  AOI22S U22342 ( .A1(n15948), .A2(gray_img[1878]), .B1(n17709), .B2(
        gray_img[590]), .O(n16511) );
  ND3S U22343 ( .I1(n16513), .I2(n16512), .I3(n16511), .O(n16514) );
  AN4B1S U22344 ( .I1(n16517), .I2(n16516), .I3(n16515), .B1(n16514), .O(
        n16542) );
  AOI22S U22345 ( .A1(n17778), .A2(gray_img[462]), .B1(n15895), .B2(
        gray_img[1502]), .O(n16522) );
  AOI22S U22346 ( .A1(n15877), .A2(gray_img[334]), .B1(n15899), .B2(
        gray_img[718]), .O(n16521) );
  AOI22S U22347 ( .A1(n15876), .A2(gray_img[1750]), .B1(n16188), .B2(
        gray_img[1246]), .O(n16520) );
  INV1S U22348 ( .I(gray_img[78]), .O(n23599) );
  MOAI1S U22349 ( .A1(n16002), .A2(n23599), .B1(n17780), .B2(gray_img[350]), 
        .O(n16519) );
  AN4B1S U22350 ( .I1(n16522), .I2(n16521), .I3(n16520), .B1(n16519), .O(
        n16540) );
  AOI22S U22351 ( .A1(n15872), .A2(gray_img[1118]), .B1(n17785), .B2(
        gray_img[1230]), .O(n16526) );
  AOI22S U22352 ( .A1(n15878), .A2(gray_img[1366]), .B1(n17787), .B2(
        gray_img[206]), .O(n16525) );
  AOI22S U22353 ( .A1(n17137), .A2(gray_img[86]), .B1(n15949), .B2(
        gray_img[1494]), .O(n16524) );
  INV1S U22354 ( .I(gray_img[1998]), .O(n23571) );
  MOAI1S U22355 ( .A1(n15894), .A2(n23571), .B1(n17786), .B2(gray_img[734]), 
        .O(n16523) );
  AN4B1S U22356 ( .I1(n16526), .I2(n16525), .I3(n16524), .B1(n16523), .O(
        n16539) );
  AOI22S U22357 ( .A1(gray_img[2006]), .A2(n15897), .B1(n17797), .B2(
        gray_img[1486]), .O(n16530) );
  AOI22S U22358 ( .A1(n17605), .A2(gray_img[1110]), .B1(n15879), .B2(
        gray_img[990]), .O(n16529) );
  AOI22S U22359 ( .A1(n17606), .A2(gray_img[342]), .B1(n15950), .B2(
        gray_img[214]), .O(n16528) );
  INV1S U22360 ( .I(gray_img[974]), .O(n22980) );
  MOAI1S U22361 ( .A1(n17718), .A2(n22980), .B1(n17796), .B2(gray_img[1358]), 
        .O(n16527) );
  AN4B1S U22362 ( .I1(n16530), .I2(n16529), .I3(n16528), .B1(n16527), .O(
        n16538) );
  MOAI1S U22363 ( .A1(n15868), .A2(n21141), .B1(n16001), .B2(gray_img[726]), 
        .O(n16533) );
  INV1S U22364 ( .I(n16531), .O(n17660) );
  INV1S U22365 ( .I(gray_img[1374]), .O(n28370) );
  MOAI1S U22366 ( .A1(n17660), .A2(n28370), .B1(n15874), .B2(gray_img[1102]), 
        .O(n16532) );
  NR2 U22367 ( .I1(n16533), .I2(n16532), .O(n16536) );
  AOI22S U22368 ( .A1(n17807), .A2(gray_img[982]), .B1(n15951), .B2(
        gray_img[1238]), .O(n16535) );
  AOI22S U22369 ( .A1(n17806), .A2(gray_img[222]), .B1(n17805), .B2(
        gray_img[1742]), .O(n16534) );
  ND3S U22370 ( .I1(n16536), .I2(n16535), .I3(n16534), .O(n16537) );
  AN4B1S U22371 ( .I1(n16540), .I2(n16539), .I3(n16538), .B1(n16537), .O(
        n16541) );
  ND2S U22372 ( .I1(n16542), .I2(n16541), .O(n16588) );
  AOI22S U22373 ( .A1(n16116), .A2(gray_img[510]), .B1(n15914), .B2(
        gray_img[1790]), .O(n16546) );
  AOI22S U22374 ( .A1(n17703), .A2(gray_img[638]), .B1(n17767), .B2(
        gray_img[1654]), .O(n16545) );
  AOI22S U22375 ( .A1(n17079), .A2(gray_img[502]), .B1(n15873), .B2(
        gray_img[2046]), .O(n16544) );
  INV1S U22376 ( .I(gray_img[886]), .O(n26385) );
  MOAI1S U22377 ( .A1(n17766), .A2(n26385), .B1(n17765), .B2(gray_img[1902]), 
        .O(n16543) );
  AN4B1S U22378 ( .I1(n16546), .I2(n16545), .I3(n16544), .B1(n16543), .O(
        n16563) );
  AOI22S U22379 ( .A1(n15898), .A2(gray_img[894]), .B1(n15911), .B2(
        gray_img[1918]), .O(n16550) );
  AOI22S U22380 ( .A1(n16137), .A2(gray_img[878]), .B1(n17744), .B2(
        gray_img[630]), .O(n16549) );
  AOI22S U22381 ( .A1(n15948), .A2(gray_img[1910]), .B1(n17709), .B2(
        gray_img[622]), .O(n16548) );
  INV1S U22382 ( .I(gray_img[1646]), .O(n25790) );
  MOAI1S U22383 ( .A1(n17381), .A2(n25790), .B1(n15908), .B2(gray_img[1662]), 
        .O(n16547) );
  AN4B1S U22384 ( .I1(n16550), .I2(n16549), .I3(n16548), .B1(n16547), .O(
        n16562) );
  AOI22S U22385 ( .A1(n15913), .A2(gray_img[1510]), .B1(n17750), .B2(
        gray_img[486]), .O(n16554) );
  AOI22S U22386 ( .A1(n16000), .A2(gray_img[1126]), .B1(n17751), .B2(
        gray_img[1638]), .O(n16553) );
  AOI22S U22387 ( .A1(n15909), .A2(gray_img[230]), .B1(gray_img[1382]), .B2(
        n15903), .O(n16552) );
  INV1S U22388 ( .I(gray_img[2022]), .O(n25846) );
  MOAI1S U22389 ( .A1(n17753), .A2(n25846), .B1(n17752), .B2(gray_img[358]), 
        .O(n16551) );
  AN4B1S U22390 ( .I1(n16554), .I2(n16553), .I3(n16552), .B1(n16551), .O(
        n16561) );
  INV1S U22391 ( .I(gray_img[614]), .O(n26200) );
  MOAI1S U22392 ( .A1(n17640), .A2(n26200), .B1(n17758), .B2(gray_img[870]), 
        .O(n16556) );
  INV1S U22393 ( .I(gray_img[1254]), .O(n28041) );
  MOAI1S U22394 ( .A1(n17518), .A2(n28041), .B1(n15901), .B2(gray_img[1894]), 
        .O(n16555) );
  NR2 U22395 ( .I1(n16556), .I2(n16555), .O(n16559) );
  AOI22S U22396 ( .A1(n15900), .A2(gray_img[998]), .B1(n17639), .B2(
        gray_img[742]), .O(n16558) );
  AOI22S U22397 ( .A1(n15902), .A2(gray_img[1766]), .B1(n15912), .B2(
        gray_img[102]), .O(n16557) );
  ND3S U22398 ( .I1(n16559), .I2(n16558), .I3(n16557), .O(n16560) );
  AOI22S U22399 ( .A1(n15872), .A2(gray_img[1150]), .B1(n17785), .B2(
        gray_img[1262]), .O(n16567) );
  AOI22S U22400 ( .A1(n15878), .A2(gray_img[1398]), .B1(n17787), .B2(
        gray_img[238]), .O(n16566) );
  AOI22S U22401 ( .A1(n17137), .A2(gray_img[118]), .B1(n15949), .B2(
        gray_img[1526]), .O(n16565) );
  INV1S U22402 ( .I(gray_img[2030]), .O(n25858) );
  MOAI1S U22403 ( .A1(n15894), .A2(n25858), .B1(n17786), .B2(gray_img[766]), 
        .O(n16564) );
  AN4B1S U22404 ( .I1(n16567), .I2(n16566), .I3(n16565), .B1(n16564), .O(
        n16573) );
  AOI22S U22405 ( .A1(n15876), .A2(gray_img[1782]), .B1(n16188), .B2(
        gray_img[1278]), .O(n16572) );
  AOI22S U22406 ( .A1(n17778), .A2(gray_img[494]), .B1(n15895), .B2(
        gray_img[1534]), .O(n16571) );
  AOI22S U22407 ( .A1(n17591), .A2(gray_img[382]), .B1(gray_img[110]), .B2(
        n17779), .O(n16569) );
  AOI22S U22408 ( .A1(n15877), .A2(gray_img[366]), .B1(n16368), .B2(
        gray_img[750]), .O(n16568) );
  ND2S U22409 ( .I1(n16569), .I2(n16568), .O(n16570) );
  AN4B1S U22410 ( .I1(n16573), .I2(n16572), .I3(n16571), .B1(n16570), .O(
        n16585) );
  AOI22S U22411 ( .A1(n15874), .A2(gray_img[1134]), .B1(n17148), .B2(
        gray_img[1406]), .O(n16577) );
  AOI22S U22412 ( .A1(n16001), .A2(gray_img[758]), .B1(n15875), .B2(
        gray_img[126]), .O(n16576) );
  AOI22S U22413 ( .A1(n17807), .A2(gray_img[1014]), .B1(n15951), .B2(
        gray_img[1270]), .O(n16575) );
  INV1S U22414 ( .I(gray_img[254]), .O(n27566) );
  MOAI1S U22415 ( .A1(n17533), .A2(n27566), .B1(n17805), .B2(gray_img[1774]), 
        .O(n16574) );
  AN4B1S U22416 ( .I1(n16577), .I2(n16576), .I3(n16575), .B1(n16574), .O(
        n16583) );
  AOI22S U22417 ( .A1(n17796), .A2(gray_img[1390]), .B1(n17795), .B2(
        gray_img[1006]), .O(n16582) );
  AOI22S U22418 ( .A1(n15897), .A2(gray_img[2038]), .B1(n17797), .B2(
        gray_img[1518]), .O(n16581) );
  AOI22S U22419 ( .A1(n17605), .A2(gray_img[1142]), .B1(n15879), .B2(
        gray_img[1022]), .O(n16579) );
  AOI22S U22420 ( .A1(n17606), .A2(gray_img[374]), .B1(n15950), .B2(
        gray_img[246]), .O(n16578) );
  ND2S U22421 ( .I1(n16579), .I2(n16578), .O(n16580) );
  AN4B1S U22422 ( .I1(n16583), .I2(n16582), .I3(n16581), .B1(n16580), .O(
        n16584) );
  ND3S U22423 ( .I1(n16586), .I2(n16585), .I3(n16584), .O(n16587) );
  AOI22S U22424 ( .A1(n16588), .A2(n17690), .B1(n17819), .B2(n16587), .O(
        n16589) );
  NR2 U22425 ( .I1(n15993), .I2(n15871), .O(n17364) );
  NR2 U22426 ( .I1(n15993), .I2(n17973), .O(n17171) );
  AOI22S U22427 ( .A1(n17584), .A2(template_reg[68]), .B1(n17583), .B2(
        template_reg[60]), .O(n16593) );
  ND2S U22428 ( .I1(n17585), .I2(template_reg[52]), .O(n16592) );
  NR2 U22429 ( .I1(n15994), .I2(n15871), .O(n17170) );
  AOI22S U22430 ( .A1(n17584), .A2(template_reg[71]), .B1(n17583), .B2(
        template_reg[63]), .O(n16599) );
  ND2S U22431 ( .I1(n17585), .I2(template_reg[55]), .O(n16598) );
  AOI22S U22432 ( .A1(n15908), .A2(gray_img[1563]), .B1(n17743), .B2(
        gray_img[1547]), .O(n16606) );
  AOI22S U22433 ( .A1(n15898), .A2(gray_img[795]), .B1(n15911), .B2(
        gray_img[1819]), .O(n16605) );
  AOI22S U22434 ( .A1(n15948), .A2(gray_img[1811]), .B1(n17709), .B2(
        gray_img[523]), .O(n16604) );
  INV1S U22435 ( .I(gray_img[531]), .O(n29054) );
  MOAI1S U22436 ( .A1(n17505), .A2(n29054), .B1(n16137), .B2(gray_img[779]), 
        .O(n16603) );
  AN4B1S U22437 ( .I1(n16606), .I2(n16605), .I3(n16604), .B1(n16603), .O(
        n16623) );
  AOI22S U22438 ( .A1(n16116), .A2(gray_img[411]), .B1(n15914), .B2(
        gray_img[1691]), .O(n16610) );
  AOI22S U22439 ( .A1(n17079), .A2(gray_img[403]), .B1(n15873), .B2(
        gray_img[1947]), .O(n16609) );
  AOI22S U22440 ( .A1(n15917), .A2(gray_img[787]), .B1(n17765), .B2(
        gray_img[1803]), .O(n16608) );
  INV1S U22441 ( .I(gray_img[539]), .O(n29068) );
  MOAI1S U22442 ( .A1(n17674), .A2(n29068), .B1(n17767), .B2(gray_img[1555]), 
        .O(n16607) );
  AN4B1S U22443 ( .I1(n16610), .I2(n16609), .I3(n16608), .B1(n16607), .O(
        n16622) );
  AOI22S U22444 ( .A1(n17752), .A2(gray_img[259]), .B1(n17696), .B2(
        gray_img[1923]), .O(n16614) );
  AOI22S U22445 ( .A1(n15913), .A2(gray_img[1411]), .B1(n17750), .B2(
        gray_img[387]), .O(n16613) );
  AOI22S U22446 ( .A1(n15909), .A2(gray_img[131]), .B1(n15903), .B2(
        gray_img[1283]), .O(n16612) );
  INV1S U22447 ( .I(gray_img[1539]), .O(n26592) );
  MOAI1S U22448 ( .A1(n15942), .A2(n26592), .B1(n16000), .B2(gray_img[1027]), 
        .O(n16611) );
  AN4B1S U22449 ( .I1(n16614), .I2(n16613), .I3(n16612), .B1(n16611), .O(
        n16621) );
  INV1S U22450 ( .I(gray_img[515]), .O(n29921) );
  MOAI1S U22451 ( .A1(n17640), .A2(n29921), .B1(n17758), .B2(gray_img[771]), 
        .O(n16616) );
  INV1S U22452 ( .I(gray_img[1155]), .O(n26631) );
  MOAI1S U22453 ( .A1(n17518), .A2(n26631), .B1(n15901), .B2(gray_img[1795]), 
        .O(n16615) );
  NR2 U22454 ( .I1(n16616), .I2(n16615), .O(n16619) );
  AOI22S U22455 ( .A1(n15900), .A2(gray_img[899]), .B1(n17639), .B2(
        gray_img[643]), .O(n16618) );
  AOI22S U22456 ( .A1(n15902), .A2(gray_img[1667]), .B1(n17478), .B2(
        gray_img[3]), .O(n16617) );
  ND3S U22457 ( .I1(n16619), .I2(n16618), .I3(n16617), .O(n16620) );
  AN4B1S U22458 ( .I1(n16623), .I2(n16622), .I3(n16621), .B1(n16620), .O(
        n16646) );
  AOI22S U22459 ( .A1(n17778), .A2(gray_img[395]), .B1(n15895), .B2(
        gray_img[1435]), .O(n16627) );
  AOI22S U22460 ( .A1(n15877), .A2(gray_img[267]), .B1(n15899), .B2(
        gray_img[651]), .O(n16626) );
  AOI22S U22461 ( .A1(n15876), .A2(gray_img[1683]), .B1(n16188), .B2(
        gray_img[1179]), .O(n16625) );
  INV1S U22462 ( .I(gray_img[11]), .O(n23422) );
  MOAI1S U22463 ( .A1(n16002), .A2(n23422), .B1(n17591), .B2(gray_img[283]), 
        .O(n16624) );
  AN4B1S U22464 ( .I1(n16627), .I2(n16626), .I3(n16625), .B1(n16624), .O(
        n16644) );
  AOI22S U22465 ( .A1(n15874), .A2(gray_img[1035]), .B1(n17148), .B2(
        gray_img[1307]), .O(n16631) );
  AOI22S U22466 ( .A1(n16001), .A2(gray_img[659]), .B1(n15896), .B2(
        gray_img[27]), .O(n16630) );
  AOI22S U22467 ( .A1(n17807), .A2(gray_img[915]), .B1(n15951), .B2(
        gray_img[1171]), .O(n16629) );
  INV1S U22468 ( .I(gray_img[155]), .O(n27868) );
  MOAI1S U22469 ( .A1(n17533), .A2(n27868), .B1(n17805), .B2(gray_img[1675]), 
        .O(n16628) );
  AN4B1S U22470 ( .I1(n16631), .I2(n16630), .I3(n16629), .B1(n16628), .O(
        n16643) );
  AOI22S U22471 ( .A1(n15897), .A2(gray_img[1939]), .B1(n17797), .B2(
        gray_img[1419]), .O(n16635) );
  AOI22S U22472 ( .A1(n17605), .A2(gray_img[1043]), .B1(n15879), .B2(
        gray_img[923]), .O(n16634) );
  AOI22S U22473 ( .A1(n17717), .A2(gray_img[275]), .B1(n15950), .B2(
        gray_img[147]), .O(n16633) );
  INV1S U22474 ( .I(gray_img[907]), .O(n29608) );
  MOAI1S U22475 ( .A1(n17718), .A2(n29608), .B1(n17796), .B2(gray_img[1291]), 
        .O(n16632) );
  AN4B1S U22476 ( .I1(n16635), .I2(n16634), .I3(n16633), .B1(n16632), .O(
        n16642) );
  INV1S U22477 ( .I(gray_img[19]), .O(n27855) );
  MOAI1S U22478 ( .A1(n15941), .A2(n27855), .B1(n15949), .B2(gray_img[1427]), 
        .O(n16637) );
  INV1S U22479 ( .I(gray_img[1299]), .O(n29751) );
  MOAI1S U22480 ( .A1(n15944), .A2(n29751), .B1(n17787), .B2(gray_img[139]), 
        .O(n16636) );
  NR2 U22481 ( .I1(n16637), .I2(n16636), .O(n16640) );
  AOI22S U22482 ( .A1(n15872), .A2(gray_img[1051]), .B1(n17785), .B2(
        gray_img[1163]), .O(n16639) );
  AOI22S U22483 ( .A1(n17786), .A2(gray_img[667]), .B1(n15866), .B2(
        gray_img[1931]), .O(n16638) );
  ND3S U22484 ( .I1(n16640), .I2(n16639), .I3(n16638), .O(n16641) );
  AN4B1S U22485 ( .I1(n16644), .I2(n16643), .I3(n16642), .B1(n16641), .O(
        n16645) );
  ND2S U22486 ( .I1(n16646), .I2(n16645), .O(n16693) );
  AOI22S U22487 ( .A1(n15908), .A2(gray_img[1595]), .B1(n17743), .B2(
        gray_img[1579]), .O(n16650) );
  AOI22S U22488 ( .A1(n15898), .A2(gray_img[827]), .B1(n15911), .B2(
        gray_img[1851]), .O(n16649) );
  AOI22S U22489 ( .A1(n16137), .A2(gray_img[811]), .B1(n17744), .B2(
        gray_img[563]), .O(n16648) );
  INV1S U22490 ( .I(gray_img[555]), .O(n28611) );
  MOAI1S U22491 ( .A1(n17745), .A2(n28611), .B1(n15948), .B2(gray_img[1843]), 
        .O(n16647) );
  AN4B1S U22492 ( .I1(n16650), .I2(n16649), .I3(n16648), .B1(n16647), .O(
        n16667) );
  AOI22S U22493 ( .A1(n16116), .A2(gray_img[443]), .B1(n15914), .B2(
        gray_img[1723]), .O(n16654) );
  AOI22S U22494 ( .A1(n17079), .A2(gray_img[435]), .B1(n15873), .B2(
        gray_img[1979]), .O(n16653) );
  AOI22S U22495 ( .A1(n15917), .A2(gray_img[819]), .B1(n17765), .B2(
        gray_img[1835]), .O(n16652) );
  INV1S U22496 ( .I(gray_img[571]), .O(n28147) );
  MOAI1S U22497 ( .A1(n17674), .A2(n28147), .B1(n17767), .B2(gray_img[1587]), 
        .O(n16651) );
  AN4B1S U22498 ( .I1(n16654), .I2(n16653), .I3(n16652), .B1(n16651), .O(
        n16666) );
  AOI22S U22499 ( .A1(n15913), .A2(gray_img[1443]), .B1(n17750), .B2(
        gray_img[419]), .O(n16658) );
  AOI22S U22500 ( .A1(n16000), .A2(gray_img[1059]), .B1(n17751), .B2(
        gray_img[1571]), .O(n16657) );
  AOI22S U22501 ( .A1(n15909), .A2(gray_img[163]), .B1(n15903), .B2(
        gray_img[1315]), .O(n16656) );
  INV1S U22502 ( .I(gray_img[1955]), .O(n26660) );
  MOAI1S U22503 ( .A1(n17753), .A2(n26660), .B1(n17752), .B2(gray_img[291]), 
        .O(n16655) );
  AN4B1S U22504 ( .I1(n16658), .I2(n16657), .I3(n16656), .B1(n16655), .O(
        n16665) );
  INV1S U22505 ( .I(gray_img[547]), .O(n28624) );
  MOAI1S U22506 ( .A1(n17640), .A2(n28624), .B1(n17758), .B2(gray_img[803]), 
        .O(n16660) );
  INV1S U22507 ( .I(gray_img[1187]), .O(n23012) );
  MOAI1S U22508 ( .A1(n17518), .A2(n23012), .B1(n15901), .B2(gray_img[1827]), 
        .O(n16659) );
  NR2 U22509 ( .I1(n16660), .I2(n16659), .O(n16663) );
  AOI22S U22510 ( .A1(n15900), .A2(gray_img[931]), .B1(n17639), .B2(
        gray_img[675]), .O(n16662) );
  AOI22S U22511 ( .A1(n15902), .A2(gray_img[1699]), .B1(n15912), .B2(
        gray_img[35]), .O(n16661) );
  ND3S U22512 ( .I1(n16663), .I2(n16662), .I3(n16661), .O(n16664) );
  AN4B1S U22513 ( .I1(n16667), .I2(n16666), .I3(n16665), .B1(n16664), .O(
        n16691) );
  AOI22S U22514 ( .A1(n15874), .A2(gray_img[1067]), .B1(n17804), .B2(
        gray_img[1339]), .O(n16672) );
  AOI22S U22515 ( .A1(n17806), .A2(gray_img[187]), .B1(n17805), .B2(
        gray_img[1707]), .O(n16671) );
  AOI22S U22516 ( .A1(n17807), .A2(gray_img[947]), .B1(n15951), .B2(
        gray_img[1203]), .O(n16670) );
  INV1S U22517 ( .I(gray_img[59]), .O(n27713) );
  MOAI1S U22518 ( .A1(n15868), .A2(n27713), .B1(n16001), .B2(gray_img[691]), 
        .O(n16669) );
  AN4B1S U22519 ( .I1(n16672), .I2(n16671), .I3(n16670), .B1(n16669), .O(
        n16689) );
  AOI22S U22520 ( .A1(n15872), .A2(gray_img[1083]), .B1(n17785), .B2(
        gray_img[1195]), .O(n16676) );
  AOI22S U22521 ( .A1(n15878), .A2(gray_img[1331]), .B1(n17787), .B2(
        gray_img[171]), .O(n16675) );
  INV2 U22522 ( .I(n15941), .O(n17329) );
  AOI22S U22523 ( .A1(n17329), .A2(gray_img[51]), .B1(n15949), .B2(
        gray_img[1459]), .O(n16674) );
  INV1S U22524 ( .I(gray_img[1963]), .O(n26673) );
  MOAI1S U22525 ( .A1(n15894), .A2(n26673), .B1(n17786), .B2(gray_img[699]), 
        .O(n16673) );
  AN4B1S U22526 ( .I1(n16676), .I2(n16675), .I3(n16674), .B1(n16673), .O(
        n16688) );
  AOI22S U22527 ( .A1(n15897), .A2(gray_img[1971]), .B1(n17797), .B2(
        gray_img[1451]), .O(n16680) );
  AOI22S U22528 ( .A1(n17605), .A2(gray_img[1075]), .B1(n15879), .B2(
        gray_img[955]), .O(n16679) );
  AOI22S U22529 ( .A1(n17717), .A2(gray_img[307]), .B1(n15950), .B2(
        gray_img[179]), .O(n16678) );
  INV1S U22530 ( .I(gray_img[939]), .O(n23212) );
  MOAI1S U22531 ( .A1(n17718), .A2(n23212), .B1(n17796), .B2(gray_img[1323]), 
        .O(n16677) );
  AN4B1S U22532 ( .I1(n16680), .I2(n16679), .I3(n16678), .B1(n16677), .O(
        n16687) );
  INV1S U22533 ( .I(gray_img[43]), .O(n26960) );
  MOAI1S U22534 ( .A1(n16002), .A2(n26960), .B1(n17780), .B2(gray_img[315]), 
        .O(n16682) );
  INV1S U22535 ( .I(gray_img[299]), .O(n27279) );
  MOAI1S U22536 ( .A1(n16518), .A2(n27279), .B1(n15899), .B2(gray_img[683]), 
        .O(n16681) );
  NR2 U22537 ( .I1(n16682), .I2(n16681), .O(n16685) );
  AOI22S U22538 ( .A1(n15876), .A2(gray_img[1715]), .B1(n16188), .B2(
        gray_img[1211]), .O(n16684) );
  AOI22S U22539 ( .A1(n17778), .A2(gray_img[427]), .B1(n15895), .B2(
        gray_img[1467]), .O(n16683) );
  ND3S U22540 ( .I1(n16685), .I2(n16684), .I3(n16683), .O(n16686) );
  AN4B1S U22541 ( .I1(n16689), .I2(n16688), .I3(n16687), .B1(n16686), .O(
        n16690) );
  ND2S U22542 ( .I1(n16691), .I2(n16690), .O(n16692) );
  AOI22S U22543 ( .A1(n16693), .A2(n17688), .B1(n17817), .B2(n16692), .O(
        n16785) );
  AOI22S U22544 ( .A1(n16116), .A2(gray_img[507]), .B1(n15914), .B2(
        gray_img[1787]), .O(n16697) );
  AOI22S U22545 ( .A1(n17703), .A2(gray_img[635]), .B1(n17767), .B2(
        gray_img[1651]), .O(n16696) );
  AOI22S U22546 ( .A1(n17079), .A2(gray_img[499]), .B1(n15873), .B2(
        gray_img[2043]), .O(n16695) );
  INV1S U22547 ( .I(gray_img[883]), .O(n26379) );
  MOAI1S U22548 ( .A1(n17766), .A2(n26379), .B1(n17765), .B2(gray_img[1899]), 
        .O(n16694) );
  AN4B1S U22549 ( .I1(n16697), .I2(n16696), .I3(n16695), .B1(n16694), .O(
        n16714) );
  AOI22S U22550 ( .A1(n15913), .A2(gray_img[1507]), .B1(n17750), .B2(
        gray_img[483]), .O(n16701) );
  AOI22S U22551 ( .A1(n16000), .A2(gray_img[1123]), .B1(n17751), .B2(
        gray_img[1635]), .O(n16700) );
  AOI22S U22552 ( .A1(n15909), .A2(gray_img[227]), .B1(n15903), .B2(
        gray_img[1379]), .O(n16699) );
  INV1S U22553 ( .I(gray_img[2019]), .O(n25840) );
  MOAI1S U22554 ( .A1(n17753), .A2(n25840), .B1(n17752), .B2(gray_img[355]), 
        .O(n16698) );
  AN4B1S U22555 ( .I1(n16701), .I2(n16700), .I3(n16699), .B1(n16698), .O(
        n16713) );
  AOI22S U22556 ( .A1(n15902), .A2(gray_img[1763]), .B1(n17478), .B2(
        gray_img[99]), .O(n16705) );
  AOI22S U22557 ( .A1(n17758), .A2(gray_img[867]), .B1(n16165), .B2(
        gray_img[611]), .O(n16704) );
  AOI22S U22558 ( .A1(n17759), .A2(gray_img[1251]), .B1(n15901), .B2(
        gray_img[1891]), .O(n16703) );
  INV1S U22559 ( .I(gray_img[739]), .O(n26166) );
  MOAI1S U22560 ( .A1(n17760), .A2(n26166), .B1(n15900), .B2(gray_img[995]), 
        .O(n16702) );
  AN4B1S U22561 ( .I1(n16705), .I2(n16704), .I3(n16703), .B1(n16702), .O(
        n16712) );
  INV1S U22562 ( .I(gray_img[891]), .O(n26392) );
  MOAI1S U22563 ( .A1(n15946), .A2(n26392), .B1(n15911), .B2(gray_img[1915]), 
        .O(n16707) );
  INV1S U22564 ( .I(gray_img[619]), .O(n26187) );
  MOAI1S U22565 ( .A1(n17745), .A2(n26187), .B1(n15948), .B2(gray_img[1907]), 
        .O(n16706) );
  NR2 U22566 ( .I1(n16707), .I2(n16706), .O(n16710) );
  AOI22S U22567 ( .A1(n15908), .A2(gray_img[1659]), .B1(n17743), .B2(
        gray_img[1643]), .O(n16709) );
  AOI22S U22568 ( .A1(n16137), .A2(gray_img[875]), .B1(n17744), .B2(
        gray_img[627]), .O(n16708) );
  ND3S U22569 ( .I1(n16710), .I2(n16709), .I3(n16708), .O(n16711) );
  AN4B1S U22570 ( .I1(n16714), .I2(n16713), .I3(n16712), .B1(n16711), .O(
        n16737) );
  AOI22S U22571 ( .A1(n15872), .A2(gray_img[1147]), .B1(n17785), .B2(
        gray_img[1259]), .O(n16718) );
  AOI22S U22572 ( .A1(n15878), .A2(gray_img[1395]), .B1(n17787), .B2(
        gray_img[235]), .O(n16717) );
  AOI22S U22573 ( .A1(n17329), .A2(gray_img[115]), .B1(n15949), .B2(
        gray_img[1523]), .O(n16716) );
  INV1S U22574 ( .I(gray_img[2027]), .O(n25852) );
  MOAI1S U22575 ( .A1(n15894), .A2(n25852), .B1(n17786), .B2(gray_img[763]), 
        .O(n16715) );
  AN4B1S U22576 ( .I1(n16718), .I2(n16717), .I3(n16716), .B1(n16715), .O(
        n16724) );
  INV1S U22577 ( .I(gray_img[1779]), .O(n26000) );
  MOAI1S U22578 ( .A1(n15947), .A2(n26000), .B1(n16188), .B2(gray_img[1275]), 
        .O(n16720) );
  INV1S U22579 ( .I(gray_img[1531]), .O(n27896) );
  MOAI1S U22580 ( .A1(n15867), .A2(n27896), .B1(n17778), .B2(gray_img[491]), 
        .O(n16719) );
  NR2 U22581 ( .I1(n16720), .I2(n16719), .O(n16723) );
  AOI22S U22582 ( .A1(n17780), .A2(gray_img[379]), .B1(n17779), .B2(
        gray_img[107]), .O(n16722) );
  INV1S U22583 ( .I(gray_img[363]), .O(n27455) );
  MOAI1S U22584 ( .A1(n16518), .A2(n27455), .B1(n15899), .B2(gray_img[747]), 
        .O(n16721) );
  AN4B1S U22585 ( .I1(n16724), .I2(n16723), .I3(n16722), .B1(n16721), .O(
        n16736) );
  AOI22S U22586 ( .A1(n15874), .A2(gray_img[1131]), .B1(n17804), .B2(
        gray_img[1403]), .O(n16728) );
  AOI22S U22587 ( .A1(n16001), .A2(gray_img[755]), .B1(n15896), .B2(
        gray_img[123]), .O(n16727) );
  AOI22S U22588 ( .A1(n17807), .A2(gray_img[1011]), .B1(n15951), .B2(
        gray_img[1267]), .O(n16726) );
  INV1S U22589 ( .I(gray_img[251]), .O(n27560) );
  MOAI1S U22590 ( .A1(n17533), .A2(n27560), .B1(n17805), .B2(gray_img[1771]), 
        .O(n16725) );
  AN4B1S U22591 ( .I1(n16728), .I2(n16727), .I3(n16726), .B1(n16725), .O(
        n16734) );
  AOI22S U22592 ( .A1(n17796), .A2(gray_img[1387]), .B1(n17795), .B2(
        gray_img[1003]), .O(n16733) );
  AOI22S U22593 ( .A1(n15897), .A2(gray_img[2035]), .B1(n17797), .B2(
        gray_img[1515]), .O(n16732) );
  AOI22S U22594 ( .A1(n17605), .A2(gray_img[1139]), .B1(n15879), .B2(
        gray_img[1019]), .O(n16730) );
  AOI22S U22595 ( .A1(n17717), .A2(gray_img[371]), .B1(n15950), .B2(
        gray_img[243]), .O(n16729) );
  ND2S U22596 ( .I1(n16730), .I2(n16729), .O(n16731) );
  AN4B1S U22597 ( .I1(n16734), .I2(n16733), .I3(n16732), .B1(n16731), .O(
        n16735) );
  AOI22S U22598 ( .A1(n15913), .A2(gray_img[1475]), .B1(n17750), .B2(
        gray_img[451]), .O(n16741) );
  AOI22S U22599 ( .A1(n16000), .A2(gray_img[1091]), .B1(n17751), .B2(
        gray_img[1603]), .O(n16740) );
  AOI22S U22600 ( .A1(n15909), .A2(gray_img[195]), .B1(n15903), .B2(
        gray_img[1347]), .O(n16739) );
  INV1S U22601 ( .I(gray_img[1987]), .O(n23552) );
  MOAI1S U22602 ( .A1(n17753), .A2(n23552), .B1(n17752), .B2(gray_img[323]), 
        .O(n16738) );
  AN4B1S U22603 ( .I1(n16741), .I2(n16740), .I3(n16739), .B1(n16738), .O(
        n16758) );
  AOI22S U22604 ( .A1(n15902), .A2(gray_img[1731]), .B1(n15912), .B2(
        gray_img[67]), .O(n16745) );
  AOI22S U22605 ( .A1(n17758), .A2(gray_img[835]), .B1(n16165), .B2(
        gray_img[579]), .O(n16744) );
  AOI22S U22606 ( .A1(n17759), .A2(gray_img[1219]), .B1(n15901), .B2(
        gray_img[1859]), .O(n16743) );
  INV1S U22607 ( .I(gray_img[707]), .O(n27138) );
  MOAI1S U22608 ( .A1(n17760), .A2(n27138), .B1(n15900), .B2(gray_img[963]), 
        .O(n16742) );
  AN4B1S U22609 ( .I1(n16745), .I2(n16744), .I3(n16743), .B1(n16742), .O(
        n16757) );
  AOI22S U22610 ( .A1(n16116), .A2(gray_img[475]), .B1(n15914), .B2(
        gray_img[1755]), .O(n16749) );
  AOI22S U22611 ( .A1(n17770), .A2(gray_img[467]), .B1(n15873), .B2(
        gray_img[2011]), .O(n16748) );
  AOI22S U22612 ( .A1(n15917), .A2(gray_img[851]), .B1(n17765), .B2(
        gray_img[1867]), .O(n16747) );
  INV1S U22613 ( .I(gray_img[1619]), .O(n25516) );
  MOAI1S U22614 ( .A1(n17704), .A2(n25516), .B1(n17703), .B2(gray_img[603]), 
        .O(n16746) );
  AN4B1S U22615 ( .I1(n16749), .I2(n16748), .I3(n16747), .B1(n16746), .O(
        n16756) );
  INV1S U22616 ( .I(gray_img[595]), .O(n27017) );
  MOAI1S U22617 ( .A1(n17505), .A2(n27017), .B1(n16137), .B2(gray_img[843]), 
        .O(n16751) );
  INV1S U22618 ( .I(gray_img[1611]), .O(n25658) );
  MOAI1S U22619 ( .A1(n17381), .A2(n25658), .B1(n15908), .B2(gray_img[1627]), 
        .O(n16750) );
  NR2 U22620 ( .I1(n16751), .I2(n16750), .O(n16754) );
  AOI22S U22621 ( .A1(n15898), .A2(gray_img[859]), .B1(n15911), .B2(
        gray_img[1883]), .O(n16753) );
  AOI22S U22622 ( .A1(n15948), .A2(gray_img[1875]), .B1(n17709), .B2(
        gray_img[587]), .O(n16752) );
  ND3S U22623 ( .I1(n16754), .I2(n16753), .I3(n16752), .O(n16755) );
  AN4B1S U22624 ( .I1(n16758), .I2(n16757), .I3(n16756), .B1(n16755), .O(
        n16781) );
  AOI22S U22625 ( .A1(n17778), .A2(gray_img[459]), .B1(n15895), .B2(
        gray_img[1499]), .O(n16762) );
  AOI22S U22626 ( .A1(n15877), .A2(gray_img[331]), .B1(n15899), .B2(
        gray_img[715]), .O(n16761) );
  AOI22S U22627 ( .A1(n15876), .A2(gray_img[1747]), .B1(n16188), .B2(
        gray_img[1243]), .O(n16760) );
  INV1S U22628 ( .I(gray_img[75]), .O(n23593) );
  MOAI1S U22629 ( .A1(n16002), .A2(n23593), .B1(n17780), .B2(gray_img[347]), 
        .O(n16759) );
  AN4B1S U22630 ( .I1(n16762), .I2(n16761), .I3(n16760), .B1(n16759), .O(
        n16779) );
  AOI22S U22631 ( .A1(n15872), .A2(gray_img[1115]), .B1(n17785), .B2(
        gray_img[1227]), .O(n16766) );
  AOI22S U22632 ( .A1(n15878), .A2(gray_img[1363]), .B1(n17787), .B2(
        gray_img[203]), .O(n16765) );
  AOI22S U22633 ( .A1(n17329), .A2(gray_img[83]), .B1(n15949), .B2(
        gray_img[1491]), .O(n16764) );
  INV1S U22634 ( .I(gray_img[1995]), .O(n23565) );
  MOAI1S U22635 ( .A1(n15894), .A2(n23565), .B1(n17786), .B2(gray_img[731]), 
        .O(n16763) );
  AN4B1S U22636 ( .I1(n16766), .I2(n16765), .I3(n16764), .B1(n16763), .O(
        n16778) );
  AOI22S U22637 ( .A1(n15897), .A2(gray_img[2003]), .B1(n17797), .B2(
        gray_img[1483]), .O(n16770) );
  AOI22S U22638 ( .A1(n17605), .A2(gray_img[1107]), .B1(n15879), .B2(
        gray_img[987]), .O(n16769) );
  AOI22S U22639 ( .A1(n17717), .A2(gray_img[339]), .B1(n15950), .B2(
        gray_img[211]), .O(n16768) );
  INV1S U22640 ( .I(gray_img[971]), .O(n22975) );
  MOAI1S U22641 ( .A1(n17718), .A2(n22975), .B1(n17796), .B2(gray_img[1355]), 
        .O(n16767) );
  AN4B1S U22642 ( .I1(n16770), .I2(n16769), .I3(n16768), .B1(n16767), .O(
        n16777) );
  MOAI1S U22643 ( .A1(n15868), .A2(n21534), .B1(n16001), .B2(gray_img[723]), 
        .O(n16772) );
  INV1S U22644 ( .I(gray_img[1371]), .O(n28364) );
  MOAI1S U22645 ( .A1(n17660), .A2(n28364), .B1(n15874), .B2(gray_img[1099]), 
        .O(n16771) );
  NR2 U22646 ( .I1(n16772), .I2(n16771), .O(n16775) );
  AOI22S U22647 ( .A1(n17807), .A2(gray_img[979]), .B1(n15951), .B2(
        gray_img[1235]), .O(n16774) );
  AOI22S U22648 ( .A1(n17806), .A2(gray_img[219]), .B1(n17805), .B2(
        gray_img[1739]), .O(n16773) );
  ND3S U22649 ( .I1(n16775), .I2(n16774), .I3(n16773), .O(n16776) );
  AN4B1S U22650 ( .I1(n16779), .I2(n16778), .I3(n16777), .B1(n16776), .O(
        n16780) );
  ND2S U22651 ( .I1(n16781), .I2(n16780), .O(n16782) );
  AOI22S U22652 ( .A1(n16783), .A2(n17819), .B1(n17690), .B2(n16782), .O(
        n16784) );
  ND2S U22653 ( .I1(n16785), .I2(n16784), .O(n16786) );
  NR2 U22654 ( .I1(n15997), .I2(n17873), .O(n17169) );
  AOI22S U22655 ( .A1(n17584), .A2(template_reg[70]), .B1(n17583), .B2(
        template_reg[62]), .O(n16789) );
  ND2S U22656 ( .I1(n17585), .I2(template_reg[54]), .O(n16788) );
  AOI22S U22657 ( .A1(n15913), .A2(gray_img[1476]), .B1(n17750), .B2(
        gray_img[452]), .O(n16796) );
  AOI22S U22658 ( .A1(n16000), .A2(gray_img[1092]), .B1(n17751), .B2(
        gray_img[1604]), .O(n16795) );
  AOI22S U22659 ( .A1(n15909), .A2(gray_img[196]), .B1(n15903), .B2(
        gray_img[1348]), .O(n16794) );
  INV1S U22660 ( .I(gray_img[1988]), .O(n23554) );
  MOAI1S U22661 ( .A1(n17753), .A2(n23554), .B1(n17752), .B2(gray_img[324]), 
        .O(n16793) );
  AN4B1S U22662 ( .I1(n16796), .I2(n16795), .I3(n16794), .B1(n16793), .O(
        n16813) );
  AOI22S U22663 ( .A1(n15902), .A2(gray_img[1732]), .B1(n17478), .B2(
        gray_img[68]), .O(n16800) );
  AOI22S U22664 ( .A1(n17758), .A2(gray_img[836]), .B1(n16165), .B2(
        gray_img[580]), .O(n16799) );
  AOI22S U22665 ( .A1(n17759), .A2(gray_img[1220]), .B1(n15901), .B2(
        gray_img[1860]), .O(n16798) );
  INV1S U22666 ( .I(gray_img[708]), .O(n27140) );
  MOAI1S U22667 ( .A1(n17760), .A2(n27140), .B1(n15900), .B2(gray_img[964]), 
        .O(n16797) );
  AN4B1S U22668 ( .I1(n16800), .I2(n16799), .I3(n16798), .B1(n16797), .O(
        n16812) );
  AOI22S U22669 ( .A1(n16116), .A2(gray_img[476]), .B1(n15914), .B2(
        gray_img[1756]), .O(n16804) );
  AOI22S U22670 ( .A1(n17079), .A2(gray_img[468]), .B1(n15873), .B2(
        gray_img[2012]), .O(n16803) );
  AOI22S U22671 ( .A1(n15917), .A2(gray_img[852]), .B1(n17765), .B2(
        gray_img[1868]), .O(n16802) );
  INV1S U22672 ( .I(gray_img[1620]), .O(n25518) );
  MOAI1S U22673 ( .A1(n17704), .A2(n25518), .B1(n17703), .B2(gray_img[604]), 
        .O(n16801) );
  AN4B1S U22674 ( .I1(n16804), .I2(n16803), .I3(n16802), .B1(n16801), .O(
        n16811) );
  INV1S U22675 ( .I(gray_img[596]), .O(n27019) );
  MOAI1S U22676 ( .A1(n17505), .A2(n27019), .B1(n16137), .B2(gray_img[844]), 
        .O(n16806) );
  INV1S U22677 ( .I(gray_img[1612]), .O(n25660) );
  MOAI1S U22678 ( .A1(n17381), .A2(n25660), .B1(n15908), .B2(gray_img[1628]), 
        .O(n16805) );
  NR2 U22679 ( .I1(n16806), .I2(n16805), .O(n16809) );
  AOI22S U22680 ( .A1(n15898), .A2(gray_img[860]), .B1(n15911), .B2(
        gray_img[1884]), .O(n16808) );
  AOI22S U22681 ( .A1(n15948), .A2(gray_img[1876]), .B1(n17709), .B2(
        gray_img[588]), .O(n16807) );
  ND3S U22682 ( .I1(n16809), .I2(n16808), .I3(n16807), .O(n16810) );
  AN4B1S U22683 ( .I1(n16813), .I2(n16812), .I3(n16811), .B1(n16810), .O(
        n16836) );
  AOI22S U22684 ( .A1(n15872), .A2(gray_img[1116]), .B1(n17785), .B2(
        gray_img[1228]), .O(n16817) );
  AOI22S U22685 ( .A1(n15878), .A2(gray_img[1364]), .B1(n17787), .B2(
        gray_img[204]), .O(n16816) );
  AOI22S U22686 ( .A1(n17329), .A2(gray_img[84]), .B1(n15949), .B2(
        gray_img[1492]), .O(n16815) );
  INV1S U22687 ( .I(gray_img[1996]), .O(n23567) );
  MOAI1S U22688 ( .A1(n15894), .A2(n23567), .B1(n17786), .B2(gray_img[732]), 
        .O(n16814) );
  AN4B1S U22689 ( .I1(n16817), .I2(n16816), .I3(n16815), .B1(n16814), .O(
        n16823) );
  AOI22S U22690 ( .A1(n15876), .A2(gray_img[1748]), .B1(n16188), .B2(
        gray_img[1244]), .O(n16822) );
  AOI22S U22691 ( .A1(n17778), .A2(gray_img[460]), .B1(n15895), .B2(
        gray_img[1500]), .O(n16821) );
  AOI22S U22692 ( .A1(n17780), .A2(gray_img[348]), .B1(n17779), .B2(
        gray_img[76]), .O(n16819) );
  AOI22S U22693 ( .A1(n15877), .A2(gray_img[332]), .B1(n15899), .B2(
        gray_img[716]), .O(n16818) );
  ND2S U22694 ( .I1(n16819), .I2(n16818), .O(n16820) );
  AN4B1S U22695 ( .I1(n16823), .I2(n16822), .I3(n16821), .B1(n16820), .O(
        n16835) );
  AOI22S U22696 ( .A1(n15897), .A2(gray_img[2004]), .B1(n17797), .B2(
        gray_img[1484]), .O(n16827) );
  AOI22S U22697 ( .A1(n17605), .A2(gray_img[1108]), .B1(n15879), .B2(
        gray_img[988]), .O(n16826) );
  AOI22S U22698 ( .A1(n17606), .A2(gray_img[340]), .B1(n15950), .B2(
        gray_img[212]), .O(n16825) );
  INV1S U22699 ( .I(gray_img[972]), .O(n22977) );
  MOAI1S U22700 ( .A1(n17718), .A2(n22977), .B1(n17796), .B2(gray_img[1356]), 
        .O(n16824) );
  AN4B1S U22701 ( .I1(n16827), .I2(n16826), .I3(n16825), .B1(n16824), .O(
        n16833) );
  AOI22S U22702 ( .A1(n16001), .A2(gray_img[724]), .B1(n15875), .B2(
        gray_img[92]), .O(n16832) );
  AOI22S U22703 ( .A1(n15874), .A2(gray_img[1100]), .B1(n17148), .B2(
        gray_img[1372]), .O(n16831) );
  AOI22S U22704 ( .A1(n17806), .A2(gray_img[220]), .B1(n17805), .B2(
        gray_img[1740]), .O(n16829) );
  AOI22S U22705 ( .A1(n17807), .A2(gray_img[980]), .B1(n15951), .B2(
        gray_img[1236]), .O(n16828) );
  ND2S U22706 ( .I1(n16829), .I2(n16828), .O(n16830) );
  AN4B1S U22707 ( .I1(n16833), .I2(n16832), .I3(n16831), .B1(n16830), .O(
        n16834) );
  ND3S U22708 ( .I1(n16836), .I2(n16835), .I3(n16834), .O(n16882) );
  AOI22S U22709 ( .A1(n15908), .A2(gray_img[1564]), .B1(n17743), .B2(
        gray_img[1548]), .O(n16840) );
  AOI22S U22710 ( .A1(n15898), .A2(gray_img[796]), .B1(n15911), .B2(
        gray_img[1820]), .O(n16839) );
  AOI22S U22711 ( .A1(n15948), .A2(gray_img[1812]), .B1(n17709), .B2(
        gray_img[524]), .O(n16838) );
  INV1S U22712 ( .I(gray_img[532]), .O(n29056) );
  MOAI1S U22713 ( .A1(n17505), .A2(n29056), .B1(n16137), .B2(gray_img[780]), 
        .O(n16837) );
  AN4B1S U22714 ( .I1(n16840), .I2(n16839), .I3(n16838), .B1(n16837), .O(
        n16857) );
  AOI22S U22715 ( .A1(n16116), .A2(gray_img[412]), .B1(n15914), .B2(
        gray_img[1692]), .O(n16844) );
  AOI22S U22716 ( .A1(n17703), .A2(gray_img[540]), .B1(n17767), .B2(
        gray_img[1556]), .O(n16843) );
  AOI22S U22717 ( .A1(n15917), .A2(gray_img[788]), .B1(n17765), .B2(
        gray_img[1804]), .O(n16842) );
  INV1S U22718 ( .I(gray_img[404]), .O(n28740) );
  MOAI1S U22719 ( .A1(n17221), .A2(n28740), .B1(n15873), .B2(gray_img[1948]), 
        .O(n16841) );
  AN4B1S U22720 ( .I1(n16844), .I2(n16843), .I3(n16842), .B1(n16841), .O(
        n16856) );
  AOI22S U22721 ( .A1(n17752), .A2(gray_img[260]), .B1(n17696), .B2(
        gray_img[1924]), .O(n16848) );
  AOI22S U22722 ( .A1(n15913), .A2(gray_img[1412]), .B1(n17750), .B2(
        gray_img[388]), .O(n16847) );
  AOI22S U22723 ( .A1(n15909), .A2(gray_img[132]), .B1(n15903), .B2(
        gray_img[1284]), .O(n16846) );
  INV1S U22724 ( .I(gray_img[1540]), .O(n26594) );
  MOAI1S U22725 ( .A1(n15942), .A2(n26594), .B1(n16000), .B2(gray_img[1028]), 
        .O(n16845) );
  AN4B1S U22726 ( .I1(n16848), .I2(n16847), .I3(n16846), .B1(n16845), .O(
        n16855) );
  INV1S U22727 ( .I(gray_img[516]), .O(n29923) );
  MOAI1S U22728 ( .A1(n17640), .A2(n29923), .B1(n17758), .B2(gray_img[772]), 
        .O(n16850) );
  INV1S U22729 ( .I(gray_img[1156]), .O(n26633) );
  MOAI1S U22730 ( .A1(n17518), .A2(n26633), .B1(n15901), .B2(gray_img[1796]), 
        .O(n16849) );
  NR2 U22731 ( .I1(n16850), .I2(n16849), .O(n16853) );
  AOI22S U22732 ( .A1(n15900), .A2(gray_img[900]), .B1(n17639), .B2(
        gray_img[644]), .O(n16852) );
  AOI22S U22733 ( .A1(n15902), .A2(gray_img[1668]), .B1(n15912), .B2(
        gray_img[4]), .O(n16851) );
  ND3S U22734 ( .I1(n16853), .I2(n16852), .I3(n16851), .O(n16854) );
  AN4B1S U22735 ( .I1(n16857), .I2(n16856), .I3(n16855), .B1(n16854), .O(
        n16880) );
  AOI22S U22736 ( .A1(n15872), .A2(gray_img[1052]), .B1(n17785), .B2(
        gray_img[1164]), .O(n16861) );
  AOI22S U22737 ( .A1(n15878), .A2(gray_img[1300]), .B1(n17787), .B2(
        gray_img[140]), .O(n16860) );
  AOI22S U22738 ( .A1(n17329), .A2(gray_img[20]), .B1(n15949), .B2(
        gray_img[1428]), .O(n16859) );
  INV1S U22739 ( .I(gray_img[1932]), .O(n29406) );
  MOAI1S U22740 ( .A1(n15894), .A2(n29406), .B1(n17786), .B2(gray_img[668]), 
        .O(n16858) );
  AN4B1S U22741 ( .I1(n16861), .I2(n16860), .I3(n16859), .B1(n16858), .O(
        n16867) );
  AOI22S U22742 ( .A1(n15876), .A2(gray_img[1684]), .B1(n16188), .B2(
        gray_img[1180]), .O(n16866) );
  AOI22S U22743 ( .A1(n17778), .A2(gray_img[396]), .B1(n15895), .B2(
        gray_img[1436]), .O(n16865) );
  AOI22S U22744 ( .A1(n17197), .A2(gray_img[284]), .B1(n17779), .B2(
        gray_img[12]), .O(n16863) );
  AOI22S U22745 ( .A1(n15877), .A2(gray_img[268]), .B1(n15899), .B2(
        gray_img[652]), .O(n16862) );
  ND2S U22746 ( .I1(n16863), .I2(n16862), .O(n16864) );
  AN4B1S U22747 ( .I1(n16867), .I2(n16866), .I3(n16865), .B1(n16864), .O(
        n16879) );
  AOI22S U22748 ( .A1(n15897), .A2(gray_img[1940]), .B1(n17797), .B2(
        gray_img[1420]), .O(n16871) );
  AOI22S U22749 ( .A1(n17605), .A2(gray_img[1044]), .B1(n15879), .B2(
        gray_img[924]), .O(n16870) );
  AOI22S U22750 ( .A1(n17717), .A2(gray_img[276]), .B1(n15950), .B2(
        gray_img[148]), .O(n16869) );
  INV1S U22751 ( .I(gray_img[908]), .O(n29610) );
  MOAI1S U22752 ( .A1(n17718), .A2(n29610), .B1(n17796), .B2(gray_img[1292]), 
        .O(n16868) );
  AN4B1S U22753 ( .I1(n16871), .I2(n16870), .I3(n16869), .B1(n16868), .O(
        n16877) );
  AOI22S U22754 ( .A1(n16001), .A2(gray_img[660]), .B1(n15875), .B2(
        gray_img[28]), .O(n16876) );
  AOI22S U22755 ( .A1(n15874), .A2(gray_img[1036]), .B1(n17148), .B2(
        gray_img[1308]), .O(n16875) );
  AOI22S U22756 ( .A1(n17806), .A2(gray_img[156]), .B1(n17805), .B2(
        gray_img[1676]), .O(n16873) );
  AOI22S U22757 ( .A1(n17807), .A2(gray_img[916]), .B1(n15951), .B2(
        gray_img[1172]), .O(n16872) );
  ND2S U22758 ( .I1(n16873), .I2(n16872), .O(n16874) );
  AN4B1S U22759 ( .I1(n16877), .I2(n16876), .I3(n16875), .B1(n16874), .O(
        n16878) );
  ND3S U22760 ( .I1(n16880), .I2(n16879), .I3(n16878), .O(n16881) );
  AOI22S U22761 ( .A1(n16882), .A2(n17690), .B1(n16881), .B2(n17688), .O(
        n16974) );
  AOI22S U22762 ( .A1(n15874), .A2(gray_img[1132]), .B1(n17148), .B2(
        gray_img[1404]), .O(n16886) );
  AOI22S U22763 ( .A1(n16001), .A2(gray_img[756]), .B1(n15896), .B2(
        gray_img[124]), .O(n16885) );
  AOI22S U22764 ( .A1(n17807), .A2(gray_img[1012]), .B1(n15951), .B2(
        gray_img[1268]), .O(n16884) );
  INV1S U22765 ( .I(gray_img[252]), .O(n27562) );
  MOAI1S U22766 ( .A1(n17533), .A2(n27562), .B1(n17805), .B2(gray_img[1772]), 
        .O(n16883) );
  AN4B1S U22767 ( .I1(n16886), .I2(n16885), .I3(n16884), .B1(n16883), .O(
        n16892) );
  AOI22S U22768 ( .A1(n17796), .A2(gray_img[1388]), .B1(n17795), .B2(
        gray_img[1004]), .O(n16891) );
  AOI22S U22769 ( .A1(n17716), .A2(gray_img[2036]), .B1(n17797), .B2(
        gray_img[1516]), .O(n16890) );
  AOI22S U22770 ( .A1(n17605), .A2(gray_img[1140]), .B1(n15879), .B2(
        gray_img[1020]), .O(n16888) );
  AOI22S U22771 ( .A1(n17798), .A2(gray_img[372]), .B1(n15950), .B2(
        gray_img[244]), .O(n16887) );
  ND2S U22772 ( .I1(n16888), .I2(n16887), .O(n16889) );
  AN4B1S U22773 ( .I1(n16892), .I2(n16891), .I3(n16890), .B1(n16889), .O(
        n16926) );
  AOI22S U22774 ( .A1(n15872), .A2(gray_img[1148]), .B1(n17785), .B2(
        gray_img[1260]), .O(n16896) );
  AOI22S U22775 ( .A1(n15878), .A2(gray_img[1396]), .B1(n17787), .B2(
        gray_img[236]), .O(n16895) );
  AOI22S U22776 ( .A1(n17329), .A2(gray_img[116]), .B1(n15949), .B2(
        gray_img[1524]), .O(n16894) );
  INV1S U22777 ( .I(gray_img[2028]), .O(n25854) );
  MOAI1S U22778 ( .A1(n15894), .A2(n25854), .B1(n17786), .B2(gray_img[764]), 
        .O(n16893) );
  AN4B1S U22779 ( .I1(n16896), .I2(n16895), .I3(n16894), .B1(n16893), .O(
        n16902) );
  AOI22S U22780 ( .A1(n15876), .A2(gray_img[1780]), .B1(n16188), .B2(
        gray_img[1276]), .O(n16901) );
  AOI22S U22781 ( .A1(n17778), .A2(gray_img[492]), .B1(n15895), .B2(
        gray_img[1532]), .O(n16900) );
  AOI22S U22782 ( .A1(n17591), .A2(gray_img[380]), .B1(n17779), .B2(
        gray_img[108]), .O(n16898) );
  AOI22S U22783 ( .A1(n15877), .A2(gray_img[364]), .B1(n15899), .B2(
        gray_img[748]), .O(n16897) );
  ND2S U22784 ( .I1(n16898), .I2(n16897), .O(n16899) );
  AN4B1S U22785 ( .I1(n16902), .I2(n16901), .I3(n16900), .B1(n16899), .O(
        n16925) );
  AOI22S U22786 ( .A1(n16116), .A2(gray_img[508]), .B1(n15914), .B2(
        gray_img[1788]), .O(n16906) );
  AOI22S U22787 ( .A1(n17703), .A2(gray_img[636]), .B1(n17767), .B2(
        gray_img[1652]), .O(n16905) );
  AOI22S U22788 ( .A1(n17079), .A2(gray_img[500]), .B1(n15873), .B2(
        gray_img[2044]), .O(n16904) );
  INV1S U22789 ( .I(gray_img[884]), .O(n26381) );
  MOAI1S U22790 ( .A1(n17766), .A2(n26381), .B1(n17765), .B2(gray_img[1900]), 
        .O(n16903) );
  AN4B1S U22791 ( .I1(n16906), .I2(n16905), .I3(n16904), .B1(n16903), .O(
        n16923) );
  AOI22S U22792 ( .A1(n15913), .A2(gray_img[1508]), .B1(n17750), .B2(
        gray_img[484]), .O(n16910) );
  AOI22S U22793 ( .A1(n15909), .A2(gray_img[228]), .B1(n15903), .B2(
        gray_img[1380]), .O(n16908) );
  INV1S U22794 ( .I(gray_img[2020]), .O(n25842) );
  MOAI1S U22795 ( .A1(n17753), .A2(n25842), .B1(n17752), .B2(gray_img[356]), 
        .O(n16907) );
  AN4B1S U22796 ( .I1(n16910), .I2(n16909), .I3(n16908), .B1(n16907), .O(
        n16922) );
  AOI22S U22797 ( .A1(n15902), .A2(gray_img[1764]), .B1(n17478), .B2(
        gray_img[100]), .O(n16914) );
  AOI22S U22798 ( .A1(n17758), .A2(gray_img[868]), .B1(n16165), .B2(
        gray_img[612]), .O(n16913) );
  AOI22S U22799 ( .A1(n17759), .A2(gray_img[1252]), .B1(n15901), .B2(
        gray_img[1892]), .O(n16912) );
  INV1S U22800 ( .I(gray_img[740]), .O(n26168) );
  MOAI1S U22801 ( .A1(n17760), .A2(n26168), .B1(n15900), .B2(gray_img[996]), 
        .O(n16911) );
  AN4B1S U22802 ( .I1(n16914), .I2(n16913), .I3(n16912), .B1(n16911), .O(
        n16921) );
  INV1S U22803 ( .I(gray_img[892]), .O(n26394) );
  MOAI1S U22804 ( .A1(n15946), .A2(n26394), .B1(n15911), .B2(gray_img[1916]), 
        .O(n16916) );
  INV1S U22805 ( .I(gray_img[620]), .O(n26185) );
  MOAI1S U22806 ( .A1(n17745), .A2(n26185), .B1(n15948), .B2(gray_img[1908]), 
        .O(n16915) );
  NR2 U22807 ( .I1(n16916), .I2(n16915), .O(n16919) );
  AOI22S U22808 ( .A1(n15908), .A2(gray_img[1660]), .B1(n17743), .B2(
        gray_img[1644]), .O(n16918) );
  AOI22S U22809 ( .A1(n16137), .A2(gray_img[876]), .B1(n17744), .B2(
        gray_img[628]), .O(n16917) );
  ND3S U22810 ( .I1(n16919), .I2(n16918), .I3(n16917), .O(n16920) );
  AN4B1S U22811 ( .I1(n16923), .I2(n16922), .I3(n16921), .B1(n16920), .O(
        n16924) );
  ND3S U22812 ( .I1(n16926), .I2(n16925), .I3(n16924), .O(n16972) );
  AOI22S U22813 ( .A1(n15908), .A2(gray_img[1596]), .B1(n17743), .B2(
        gray_img[1580]), .O(n16930) );
  AOI22S U22814 ( .A1(n15898), .A2(gray_img[828]), .B1(n15911), .B2(
        gray_img[1852]), .O(n16929) );
  AOI22S U22815 ( .A1(n16137), .A2(gray_img[812]), .B1(n17744), .B2(
        gray_img[564]), .O(n16928) );
  INV1S U22816 ( .I(gray_img[556]), .O(n28613) );
  MOAI1S U22817 ( .A1(n17745), .A2(n28613), .B1(n15948), .B2(gray_img[1844]), 
        .O(n16927) );
  AN4B1S U22818 ( .I1(n16930), .I2(n16929), .I3(n16928), .B1(n16927), .O(
        n16947) );
  AOI22S U22819 ( .A1(n16116), .A2(gray_img[444]), .B1(n15914), .B2(
        gray_img[1724]), .O(n16934) );
  AOI22S U22820 ( .A1(n17703), .A2(gray_img[572]), .B1(n17767), .B2(
        gray_img[1588]), .O(n16933) );
  AOI22S U22821 ( .A1(n17079), .A2(gray_img[436]), .B1(n15873), .B2(
        gray_img[1980]), .O(n16932) );
  INV1S U22822 ( .I(gray_img[820]), .O(n26104) );
  MOAI1S U22823 ( .A1(n17766), .A2(n26104), .B1(n17765), .B2(gray_img[1836]), 
        .O(n16931) );
  AN4B1S U22824 ( .I1(n16934), .I2(n16933), .I3(n16932), .B1(n16931), .O(
        n16946) );
  AOI22S U22825 ( .A1(n15913), .A2(gray_img[1444]), .B1(n17750), .B2(
        gray_img[420]), .O(n16938) );
  AOI22S U22826 ( .A1(n16000), .A2(gray_img[1060]), .B1(n17751), .B2(
        gray_img[1572]), .O(n16937) );
  AOI22S U22827 ( .A1(n15909), .A2(gray_img[164]), .B1(n15903), .B2(
        gray_img[1316]), .O(n16936) );
  INV1S U22828 ( .I(gray_img[1956]), .O(n26662) );
  MOAI1S U22829 ( .A1(n17753), .A2(n26662), .B1(n17752), .B2(gray_img[292]), 
        .O(n16935) );
  AN4B1S U22830 ( .I1(n16938), .I2(n16937), .I3(n16936), .B1(n16935), .O(
        n16945) );
  INV1S U22831 ( .I(gray_img[548]), .O(n28626) );
  MOAI1S U22832 ( .A1(n17640), .A2(n28626), .B1(n17758), .B2(gray_img[804]), 
        .O(n16940) );
  INV1S U22833 ( .I(gray_img[1188]), .O(n23014) );
  MOAI1S U22834 ( .A1(n17518), .A2(n23014), .B1(n15901), .B2(gray_img[1828]), 
        .O(n16939) );
  NR2 U22835 ( .I1(n16940), .I2(n16939), .O(n16943) );
  AOI22S U22836 ( .A1(n15900), .A2(gray_img[932]), .B1(n17639), .B2(
        gray_img[676]), .O(n16942) );
  AOI22S U22837 ( .A1(n15902), .A2(gray_img[1700]), .B1(n17478), .B2(
        gray_img[36]), .O(n16941) );
  ND3S U22838 ( .I1(n16943), .I2(n16942), .I3(n16941), .O(n16944) );
  AN4B1S U22839 ( .I1(n16947), .I2(n16946), .I3(n16945), .B1(n16944), .O(
        n16970) );
  AOI22S U22840 ( .A1(n15872), .A2(gray_img[1084]), .B1(n17785), .B2(
        gray_img[1196]), .O(n16951) );
  AOI22S U22841 ( .A1(n15878), .A2(gray_img[1332]), .B1(n17787), .B2(
        gray_img[172]), .O(n16950) );
  AOI22S U22842 ( .A1(n17329), .A2(gray_img[52]), .B1(n15949), .B2(
        gray_img[1460]), .O(n16949) );
  INV1S U22843 ( .I(gray_img[1964]), .O(n26675) );
  MOAI1S U22844 ( .A1(n15894), .A2(n26675), .B1(n17786), .B2(gray_img[700]), 
        .O(n16948) );
  AN4B1S U22845 ( .I1(n16951), .I2(n16950), .I3(n16949), .B1(n16948), .O(
        n16957) );
  AOI22S U22846 ( .A1(n15876), .A2(gray_img[1716]), .B1(n16188), .B2(
        gray_img[1212]), .O(n16956) );
  AOI22S U22847 ( .A1(n17778), .A2(gray_img[428]), .B1(n15895), .B2(
        gray_img[1468]), .O(n16955) );
  AOI22S U22848 ( .A1(n17591), .A2(gray_img[316]), .B1(n17779), .B2(
        gray_img[44]), .O(n16953) );
  AOI22S U22849 ( .A1(n15877), .A2(gray_img[300]), .B1(n15899), .B2(
        gray_img[684]), .O(n16952) );
  ND2S U22850 ( .I1(n16953), .I2(n16952), .O(n16954) );
  AN4B1S U22851 ( .I1(n16957), .I2(n16956), .I3(n16955), .B1(n16954), .O(
        n16969) );
  AOI22S U22852 ( .A1(n15897), .A2(gray_img[1972]), .B1(n17797), .B2(
        gray_img[1452]), .O(n16961) );
  AOI22S U22853 ( .A1(n17605), .A2(gray_img[1076]), .B1(n15879), .B2(
        gray_img[956]), .O(n16960) );
  AOI22S U22854 ( .A1(n17606), .A2(gray_img[308]), .B1(n15950), .B2(
        gray_img[180]), .O(n16959) );
  INV1S U22855 ( .I(gray_img[940]), .O(n23214) );
  MOAI1S U22856 ( .A1(n17718), .A2(n23214), .B1(n17796), .B2(gray_img[1324]), 
        .O(n16958) );
  AN4B1S U22857 ( .I1(n16961), .I2(n16960), .I3(n16959), .B1(n16958), .O(
        n16967) );
  AOI22S U22858 ( .A1(n16001), .A2(gray_img[692]), .B1(n15896), .B2(
        gray_img[60]), .O(n16966) );
  AOI22S U22859 ( .A1(n17723), .A2(gray_img[1068]), .B1(n17148), .B2(
        gray_img[1340]), .O(n16965) );
  AOI22S U22860 ( .A1(n17806), .A2(gray_img[188]), .B1(n17805), .B2(
        gray_img[1708]), .O(n16963) );
  AOI22S U22861 ( .A1(n17807), .A2(gray_img[948]), .B1(n15951), .B2(
        gray_img[1204]), .O(n16962) );
  ND2S U22862 ( .I1(n16963), .I2(n16962), .O(n16964) );
  AN4B1S U22863 ( .I1(n16967), .I2(n16966), .I3(n16965), .B1(n16964), .O(
        n16968) );
  ND3S U22864 ( .I1(n16970), .I2(n16969), .I3(n16968), .O(n16971) );
  AOI22S U22865 ( .A1(n16972), .A2(n17819), .B1(n16971), .B2(n17817), .O(
        n16973) );
  NR2 U22866 ( .I1(n15996), .I2(n15943), .O(n17168) );
  AOI22S U22867 ( .A1(n17584), .A2(template_reg[69]), .B1(n17583), .B2(
        template_reg[61]), .O(n16977) );
  ND2S U22868 ( .I1(n17585), .I2(template_reg[53]), .O(n16976) );
  AOI22S U22869 ( .A1(n15913), .A2(gray_img[1477]), .B1(n17750), .B2(
        gray_img[453]), .O(n16984) );
  AOI22S U22870 ( .A1(n16000), .A2(gray_img[1093]), .B1(n17751), .B2(
        gray_img[1605]), .O(n16983) );
  AOI22S U22871 ( .A1(n15909), .A2(gray_img[197]), .B1(n15903), .B2(
        gray_img[1349]), .O(n16982) );
  INV1S U22872 ( .I(gray_img[1989]), .O(n23556) );
  MOAI1S U22873 ( .A1(n17753), .A2(n23556), .B1(n17752), .B2(gray_img[325]), 
        .O(n16981) );
  AN4B1S U22874 ( .I1(n16984), .I2(n16983), .I3(n16982), .B1(n16981), .O(
        n17001) );
  AOI22S U22875 ( .A1(n15902), .A2(gray_img[1733]), .B1(n17478), .B2(
        gray_img[69]), .O(n16988) );
  AOI22S U22876 ( .A1(n17758), .A2(gray_img[837]), .B1(n16165), .B2(
        gray_img[581]), .O(n16987) );
  AOI22S U22877 ( .A1(n17759), .A2(gray_img[1221]), .B1(n15901), .B2(
        gray_img[1861]), .O(n16986) );
  INV1S U22878 ( .I(gray_img[709]), .O(n27142) );
  MOAI1S U22879 ( .A1(n17760), .A2(n27142), .B1(n15900), .B2(gray_img[965]), 
        .O(n16985) );
  AN4B1S U22880 ( .I1(n16988), .I2(n16987), .I3(n16986), .B1(n16985), .O(
        n17000) );
  AOI22S U22881 ( .A1(n16116), .A2(gray_img[477]), .B1(n15914), .B2(
        gray_img[1757]), .O(n16992) );
  AOI22S U22882 ( .A1(n17079), .A2(gray_img[469]), .B1(n15873), .B2(
        gray_img[2013]), .O(n16991) );
  AOI22S U22883 ( .A1(n15917), .A2(gray_img[853]), .B1(n17765), .B2(
        gray_img[1869]), .O(n16990) );
  INV1S U22884 ( .I(gray_img[1621]), .O(n25520) );
  MOAI1S U22885 ( .A1(n17704), .A2(n25520), .B1(n17703), .B2(gray_img[605]), 
        .O(n16989) );
  AN4B1S U22886 ( .I1(n16992), .I2(n16991), .I3(n16990), .B1(n16989), .O(
        n16999) );
  INV1S U22887 ( .I(gray_img[597]), .O(n27021) );
  MOAI1S U22888 ( .A1(n17505), .A2(n27021), .B1(n16137), .B2(gray_img[845]), 
        .O(n16994) );
  INV1S U22889 ( .I(gray_img[1613]), .O(n25662) );
  MOAI1S U22890 ( .A1(n17381), .A2(n25662), .B1(n15908), .B2(gray_img[1629]), 
        .O(n16993) );
  NR2 U22891 ( .I1(n16994), .I2(n16993), .O(n16997) );
  AOI22S U22892 ( .A1(n15898), .A2(gray_img[861]), .B1(n15911), .B2(
        gray_img[1885]), .O(n16996) );
  AOI22S U22893 ( .A1(n15948), .A2(gray_img[1877]), .B1(n17709), .B2(
        gray_img[589]), .O(n16995) );
  ND3S U22894 ( .I1(n16997), .I2(n16996), .I3(n16995), .O(n16998) );
  AN4B1S U22895 ( .I1(n17001), .I2(n17000), .I3(n16999), .B1(n16998), .O(
        n17024) );
  AOI22S U22896 ( .A1(n15872), .A2(gray_img[1117]), .B1(n17785), .B2(
        gray_img[1229]), .O(n17005) );
  AOI22S U22897 ( .A1(n15878), .A2(gray_img[1365]), .B1(n17787), .B2(
        gray_img[205]), .O(n17004) );
  AOI22S U22898 ( .A1(n17137), .A2(gray_img[85]), .B1(n15949), .B2(
        gray_img[1493]), .O(n17003) );
  INV1S U22899 ( .I(gray_img[1997]), .O(n23569) );
  MOAI1S U22900 ( .A1(n15894), .A2(n23569), .B1(n17786), .B2(gray_img[733]), 
        .O(n17002) );
  AN4B1S U22901 ( .I1(n17005), .I2(n17004), .I3(n17003), .B1(n17002), .O(
        n17011) );
  AOI22S U22902 ( .A1(n15876), .A2(gray_img[1749]), .B1(n16188), .B2(
        gray_img[1245]), .O(n17010) );
  AOI22S U22903 ( .A1(n17778), .A2(gray_img[461]), .B1(n15895), .B2(
        gray_img[1501]), .O(n17009) );
  AOI22S U22904 ( .A1(n17780), .A2(gray_img[349]), .B1(n17779), .B2(
        gray_img[77]), .O(n17007) );
  AOI22S U22905 ( .A1(n15877), .A2(gray_img[333]), .B1(n15899), .B2(
        gray_img[717]), .O(n17006) );
  ND2S U22906 ( .I1(n17007), .I2(n17006), .O(n17008) );
  AN4B1S U22907 ( .I1(n17011), .I2(n17010), .I3(n17009), .B1(n17008), .O(
        n17023) );
  AOI22S U22908 ( .A1(gray_img[2005]), .A2(n15897), .B1(n17797), .B2(
        gray_img[1485]), .O(n17015) );
  AOI22S U22909 ( .A1(n17605), .A2(gray_img[1109]), .B1(n15879), .B2(
        gray_img[989]), .O(n17014) );
  AOI22S U22910 ( .A1(n17606), .A2(gray_img[341]), .B1(n15950), .B2(
        gray_img[213]), .O(n17013) );
  INV1S U22911 ( .I(gray_img[973]), .O(n27175) );
  MOAI1S U22912 ( .A1(n17718), .A2(n27175), .B1(n17796), .B2(gray_img[1357]), 
        .O(n17012) );
  AN4B1S U22913 ( .I1(n17015), .I2(n17014), .I3(n17013), .B1(n17012), .O(
        n17021) );
  AOI22S U22914 ( .A1(n16001), .A2(gray_img[725]), .B1(n15896), .B2(
        gray_img[93]), .O(n17020) );
  AOI22S U22915 ( .A1(n17723), .A2(gray_img[1101]), .B1(n17148), .B2(
        gray_img[1373]), .O(n17019) );
  AOI22S U22916 ( .A1(n17806), .A2(gray_img[221]), .B1(n17805), .B2(
        gray_img[1741]), .O(n17017) );
  AOI22S U22917 ( .A1(n17807), .A2(gray_img[981]), .B1(n15951), .B2(
        gray_img[1237]), .O(n17016) );
  ND2S U22918 ( .I1(n17017), .I2(n17016), .O(n17018) );
  AN4B1S U22919 ( .I1(n17021), .I2(n17020), .I3(n17019), .B1(n17018), .O(
        n17022) );
  ND3S U22920 ( .I1(n17024), .I2(n17023), .I3(n17022), .O(n17070) );
  AOI22S U22921 ( .A1(n15898), .A2(gray_img[797]), .B1(n15911), .B2(
        gray_img[1821]), .O(n17028) );
  AOI22S U22922 ( .A1(n15908), .A2(gray_img[1565]), .B1(n17743), .B2(
        gray_img[1549]), .O(n17027) );
  AOI22S U22923 ( .A1(n15948), .A2(gray_img[1813]), .B1(n17709), .B2(
        gray_img[525]), .O(n17026) );
  INV1S U22924 ( .I(gray_img[533]), .O(n29058) );
  MOAI1S U22925 ( .A1(n17505), .A2(n29058), .B1(n16137), .B2(gray_img[781]), 
        .O(n17025) );
  AN4B1S U22926 ( .I1(n17028), .I2(n17027), .I3(n17026), .B1(n17025), .O(
        n17045) );
  AOI22S U22927 ( .A1(n15913), .A2(gray_img[1413]), .B1(n17750), .B2(
        gray_img[389]), .O(n17032) );
  AOI22S U22928 ( .A1(n15909), .A2(gray_img[133]), .B1(n15903), .B2(
        gray_img[1285]), .O(n17031) );
  AOI22S U22929 ( .A1(n17696), .A2(gray_img[1925]), .B1(n17752), .B2(
        gray_img[261]), .O(n17030) );
  INV1S U22930 ( .I(gray_img[1541]), .O(n26596) );
  MOAI1S U22931 ( .A1(n15942), .A2(n26596), .B1(n16000), .B2(gray_img[1029]), 
        .O(n17029) );
  AN4B1S U22932 ( .I1(n17032), .I2(n17031), .I3(n17030), .B1(n17029), .O(
        n17044) );
  AOI22S U22933 ( .A1(n16116), .A2(gray_img[413]), .B1(gray_img[1693]), .B2(
        n15914), .O(n17036) );
  AOI22S U22934 ( .A1(n15917), .A2(gray_img[789]), .B1(n17765), .B2(
        gray_img[1805]), .O(n17035) );
  AOI22S U22935 ( .A1(n17767), .A2(gray_img[1557]), .B1(n17703), .B2(
        gray_img[541]), .O(n17034) );
  INV1S U22936 ( .I(gray_img[405]), .O(n28742) );
  MOAI1S U22937 ( .A1(n17221), .A2(n28742), .B1(n15873), .B2(gray_img[1949]), 
        .O(n17033) );
  AN4B1S U22938 ( .I1(n17036), .I2(n17035), .I3(n17034), .B1(n17033), .O(
        n17043) );
  INV1S U22939 ( .I(gray_img[517]), .O(n29925) );
  MOAI1S U22940 ( .A1(n17640), .A2(n29925), .B1(n17758), .B2(gray_img[773]), 
        .O(n17038) );
  INV1S U22941 ( .I(gray_img[1797]), .O(n29395) );
  MOAI1S U22942 ( .A1(n15940), .A2(n29395), .B1(n17759), .B2(gray_img[1157]), 
        .O(n17037) );
  NR2 U22943 ( .I1(n17038), .I2(n17037), .O(n17041) );
  AOI22S U22944 ( .A1(n15900), .A2(gray_img[901]), .B1(n17639), .B2(
        gray_img[645]), .O(n17040) );
  AOI22S U22945 ( .A1(n15902), .A2(gray_img[1669]), .B1(n15912), .B2(
        gray_img[5]), .O(n17039) );
  ND3S U22946 ( .I1(n17041), .I2(n17040), .I3(n17039), .O(n17042) );
  AOI22S U22947 ( .A1(n15872), .A2(gray_img[1053]), .B1(n17785), .B2(
        gray_img[1165]), .O(n17049) );
  AOI22S U22948 ( .A1(n15878), .A2(gray_img[1301]), .B1(n17787), .B2(
        gray_img[141]), .O(n17048) );
  AOI22S U22949 ( .A1(n17137), .A2(gray_img[21]), .B1(n15949), .B2(
        gray_img[1429]), .O(n17047) );
  INV1S U22950 ( .I(gray_img[669]), .O(n29071) );
  MOAI1S U22951 ( .A1(n29071), .A2(n16003), .B1(n15866), .B2(gray_img[1933]), 
        .O(n17046) );
  AN4B1S U22952 ( .I1(n17049), .I2(n17048), .I3(n17047), .B1(n17046), .O(
        n17055) );
  AOI22S U22953 ( .A1(n15876), .A2(gray_img[1685]), .B1(n16188), .B2(
        gray_img[1181]), .O(n17054) );
  AOI22S U22954 ( .A1(n17778), .A2(gray_img[397]), .B1(n15895), .B2(
        gray_img[1437]), .O(n17053) );
  AOI22S U22955 ( .A1(n17591), .A2(gray_img[285]), .B1(n17779), .B2(
        gray_img[13]), .O(n17051) );
  AOI22S U22956 ( .A1(n15877), .A2(gray_img[269]), .B1(n16368), .B2(
        gray_img[653]), .O(n17050) );
  ND2S U22957 ( .I1(n17051), .I2(n17050), .O(n17052) );
  AN4B1S U22958 ( .I1(n17055), .I2(n17054), .I3(n17053), .B1(n17052), .O(
        n17067) );
  AOI22S U22959 ( .A1(n15897), .A2(gray_img[1941]), .B1(n17797), .B2(
        gray_img[1421]), .O(n17059) );
  AOI22S U22960 ( .A1(n17605), .A2(gray_img[1045]), .B1(n15879), .B2(
        gray_img[925]), .O(n17058) );
  AOI22S U22961 ( .A1(n17717), .A2(gray_img[277]), .B1(n15950), .B2(
        gray_img[149]), .O(n17057) );
  INV1S U22962 ( .I(gray_img[909]), .O(n29612) );
  MOAI1S U22963 ( .A1(n17718), .A2(n29612), .B1(n17796), .B2(gray_img[1293]), 
        .O(n17056) );
  AN4B1S U22964 ( .I1(n17059), .I2(n17058), .I3(n17057), .B1(n17056), .O(
        n17065) );
  AOI22S U22965 ( .A1(n16001), .A2(gray_img[661]), .B1(n15896), .B2(
        gray_img[29]), .O(n17064) );
  AOI22S U22966 ( .A1(n17723), .A2(gray_img[1037]), .B1(n17148), .B2(
        gray_img[1309]), .O(n17063) );
  AOI22S U22967 ( .A1(n17806), .A2(gray_img[157]), .B1(n17805), .B2(
        gray_img[1677]), .O(n17061) );
  AOI22S U22968 ( .A1(n17807), .A2(gray_img[917]), .B1(n15951), .B2(
        gray_img[1173]), .O(n17060) );
  ND2S U22969 ( .I1(n17061), .I2(n17060), .O(n17062) );
  AN4B1S U22970 ( .I1(n17065), .I2(n17064), .I3(n17063), .B1(n17062), .O(
        n17066) );
  ND3S U22971 ( .I1(n17068), .I2(n17067), .I3(n17066), .O(n17069) );
  AOI22S U22972 ( .A1(n17070), .A2(n17690), .B1(n17688), .B2(n17069), .O(
        n17165) );
  AOI22S U22973 ( .A1(n15898), .A2(gray_img[829]), .B1(n15911), .B2(
        gray_img[1853]), .O(n17074) );
  AOI22S U22974 ( .A1(n15908), .A2(gray_img[1597]), .B1(n17743), .B2(
        gray_img[1581]), .O(n17073) );
  INV1S U22975 ( .I(gray_img[557]), .O(n28615) );
  MOAI1S U22976 ( .A1(n17745), .A2(n28615), .B1(n15948), .B2(gray_img[1845]), 
        .O(n17071) );
  AOI22S U22977 ( .A1(n15913), .A2(gray_img[1445]), .B1(n17750), .B2(
        gray_img[421]), .O(n17078) );
  AOI22S U22978 ( .A1(n16000), .A2(gray_img[1061]), .B1(n17751), .B2(
        gray_img[1573]), .O(n17077) );
  AOI22S U22979 ( .A1(n15909), .A2(gray_img[165]), .B1(n15903), .B2(
        gray_img[1317]), .O(n17076) );
  INV1S U22980 ( .I(gray_img[293]), .O(n27271) );
  MOAI1S U22981 ( .A1(n15999), .A2(n27271), .B1(n17696), .B2(gray_img[1957]), 
        .O(n17075) );
  AN4B1S U22982 ( .I1(n17078), .I2(n17077), .I3(n17076), .B1(n17075), .O(
        n17091) );
  AOI22S U22983 ( .A1(n16116), .A2(gray_img[445]), .B1(n15914), .B2(
        gray_img[1725]), .O(n17083) );
  AOI22S U22984 ( .A1(n17079), .A2(gray_img[437]), .B1(n15873), .B2(
        gray_img[1981]), .O(n17082) );
  AOI22S U22985 ( .A1(n17767), .A2(gray_img[1589]), .B1(n17703), .B2(
        gray_img[573]), .O(n17081) );
  INV1S U22986 ( .I(gray_img[821]), .O(n26106) );
  MOAI1S U22987 ( .A1(n17766), .A2(n26106), .B1(n17765), .B2(gray_img[1837]), 
        .O(n17080) );
  INV1S U22988 ( .I(gray_img[549]), .O(n28628) );
  MOAI1S U22989 ( .A1(n17640), .A2(n28628), .B1(n17758), .B2(gray_img[805]), 
        .O(n17085) );
  INV1S U22990 ( .I(gray_img[1189]), .O(n23016) );
  MOAI1S U22991 ( .A1(n17518), .A2(n23016), .B1(n15901), .B2(gray_img[1829]), 
        .O(n17084) );
  NR2 U22992 ( .I1(n17085), .I2(n17084), .O(n17088) );
  AOI22S U22993 ( .A1(n15900), .A2(gray_img[933]), .B1(n17639), .B2(
        gray_img[677]), .O(n17087) );
  AOI22S U22994 ( .A1(n15902), .A2(gray_img[1701]), .B1(n17478), .B2(
        gray_img[37]), .O(n17086) );
  ND3S U22995 ( .I1(n17088), .I2(n17087), .I3(n17086), .O(n17089) );
  AN4B1S U22996 ( .I1(n17092), .I2(n17091), .I3(n17090), .B1(n17089), .O(
        n17115) );
  AOI22S U22997 ( .A1(n15872), .A2(gray_img[1085]), .B1(n17785), .B2(
        gray_img[1197]), .O(n17096) );
  AOI22S U22998 ( .A1(gray_img[1333]), .A2(n15878), .B1(n17787), .B2(
        gray_img[173]), .O(n17095) );
  AOI22S U22999 ( .A1(n17137), .A2(gray_img[53]), .B1(n15949), .B2(
        gray_img[1461]), .O(n17094) );
  INV1S U23000 ( .I(gray_img[1965]), .O(n26677) );
  MOAI1S U23001 ( .A1(n15894), .A2(n26677), .B1(n17786), .B2(gray_img[701]), 
        .O(n17093) );
  AN4B1S U23002 ( .I1(n17096), .I2(n17095), .I3(n17094), .B1(n17093), .O(
        n17102) );
  AOI22S U23003 ( .A1(n15876), .A2(gray_img[1717]), .B1(n16188), .B2(
        gray_img[1213]), .O(n17101) );
  AOI22S U23004 ( .A1(n17778), .A2(gray_img[429]), .B1(n15895), .B2(
        gray_img[1469]), .O(n17100) );
  AOI22S U23005 ( .A1(n17591), .A2(gray_img[317]), .B1(n17779), .B2(
        gray_img[45]), .O(n17098) );
  AOI22S U23006 ( .A1(n15877), .A2(gray_img[301]), .B1(n16368), .B2(
        gray_img[685]), .O(n17097) );
  ND2S U23007 ( .I1(n17098), .I2(n17097), .O(n17099) );
  AN4B1S U23008 ( .I1(n17102), .I2(n17101), .I3(n17100), .B1(n17099), .O(
        n17114) );
  AOI22S U23009 ( .A1(n15897), .A2(gray_img[1973]), .B1(n17797), .B2(
        gray_img[1453]), .O(n17106) );
  AOI22S U23010 ( .A1(n17605), .A2(gray_img[1077]), .B1(n15879), .B2(
        gray_img[957]), .O(n17105) );
  AOI22S U23011 ( .A1(n17606), .A2(gray_img[309]), .B1(n15950), .B2(
        gray_img[181]), .O(n17104) );
  INV1S U23012 ( .I(gray_img[941]), .O(n23216) );
  MOAI1S U23013 ( .A1(n17718), .A2(n23216), .B1(n17796), .B2(gray_img[1325]), 
        .O(n17103) );
  AN4B1S U23014 ( .I1(n17106), .I2(n17105), .I3(n17104), .B1(n17103), .O(
        n17112) );
  AOI22S U23015 ( .A1(n16001), .A2(gray_img[693]), .B1(n15896), .B2(
        gray_img[61]), .O(n17111) );
  AOI22S U23016 ( .A1(n17723), .A2(gray_img[1069]), .B1(n17148), .B2(
        gray_img[1341]), .O(n17110) );
  AOI22S U23017 ( .A1(n17806), .A2(gray_img[189]), .B1(n17805), .B2(
        gray_img[1709]), .O(n17108) );
  AOI22S U23018 ( .A1(n17807), .A2(gray_img[949]), .B1(n15951), .B2(
        gray_img[1205]), .O(n17107) );
  ND2S U23019 ( .I1(n17108), .I2(n17107), .O(n17109) );
  AN4B1S U23020 ( .I1(n17112), .I2(n17111), .I3(n17110), .B1(n17109), .O(
        n17113) );
  ND3S U23021 ( .I1(n17115), .I2(n17114), .I3(n17113), .O(n17163) );
  AOI22S U23022 ( .A1(n16116), .A2(gray_img[509]), .B1(n15914), .B2(
        gray_img[1789]), .O(n17119) );
  AOI22S U23023 ( .A1(n15917), .A2(gray_img[885]), .B1(n17765), .B2(
        gray_img[1901]), .O(n17118) );
  AOI22S U23024 ( .A1(n17767), .A2(gray_img[1653]), .B1(n17703), .B2(
        gray_img[637]), .O(n17117) );
  INV1S U23025 ( .I(gray_img[501]), .O(n27606) );
  MOAI1S U23026 ( .A1(n17221), .A2(n27606), .B1(n15873), .B2(gray_img[2045]), 
        .O(n17116) );
  AN4B1S U23027 ( .I1(n17119), .I2(n17118), .I3(n17117), .B1(n17116), .O(
        n17136) );
  AOI22S U23028 ( .A1(n15913), .A2(gray_img[1509]), .B1(n17750), .B2(
        gray_img[485]), .O(n17123) );
  AOI22S U23029 ( .A1(n16000), .A2(gray_img[1125]), .B1(n17751), .B2(
        gray_img[1637]), .O(n17122) );
  AOI22S U23030 ( .A1(n15909), .A2(gray_img[229]), .B1(gray_img[1381]), .B2(
        n15903), .O(n17121) );
  INV1S U23031 ( .I(gray_img[2021]), .O(n25844) );
  MOAI1S U23032 ( .A1(n17753), .A2(n25844), .B1(n17752), .B2(gray_img[357]), 
        .O(n17120) );
  AN4B1S U23033 ( .I1(n17123), .I2(n17122), .I3(n17121), .B1(n17120), .O(
        n17135) );
  AOI22S U23034 ( .A1(n15898), .A2(gray_img[893]), .B1(n15911), .B2(
        gray_img[1917]), .O(n17127) );
  AOI22S U23035 ( .A1(n15948), .A2(gray_img[1909]), .B1(n17709), .B2(
        gray_img[621]), .O(n17126) );
  AOI22S U23036 ( .A1(n17744), .A2(gray_img[629]), .B1(n16137), .B2(
        gray_img[877]), .O(n17125) );
  INV1S U23037 ( .I(gray_img[1645]), .O(n25788) );
  MOAI1S U23038 ( .A1(n17381), .A2(n25788), .B1(n15908), .B2(gray_img[1661]), 
        .O(n17124) );
  INV1S U23039 ( .I(gray_img[613]), .O(n26170) );
  MOAI1S U23040 ( .A1(n17640), .A2(n26170), .B1(n17758), .B2(gray_img[869]), 
        .O(n17129) );
  INV1S U23041 ( .I(gray_img[1253]), .O(n28039) );
  MOAI1S U23042 ( .A1(n17518), .A2(n28039), .B1(n15901), .B2(gray_img[1893]), 
        .O(n17128) );
  NR2 U23043 ( .I1(n17129), .I2(n17128), .O(n17132) );
  AOI22S U23044 ( .A1(n15900), .A2(gray_img[997]), .B1(n17639), .B2(
        gray_img[741]), .O(n17131) );
  AOI22S U23045 ( .A1(n15902), .A2(gray_img[1765]), .B1(n15912), .B2(
        gray_img[101]), .O(n17130) );
  ND3S U23046 ( .I1(n17132), .I2(n17131), .I3(n17130), .O(n17133) );
  AN4B1 U23047 ( .I1(n17136), .I2(n17135), .I3(n17134), .B1(n17133), .O(n17161) );
  AOI22S U23048 ( .A1(n15872), .A2(gray_img[1149]), .B1(n17785), .B2(
        gray_img[1261]), .O(n17141) );
  AOI22S U23049 ( .A1(n15878), .A2(gray_img[1397]), .B1(n17787), .B2(
        gray_img[237]), .O(n17140) );
  AOI22S U23050 ( .A1(n17137), .A2(gray_img[117]), .B1(n15949), .B2(
        gray_img[1525]), .O(n17139) );
  INV1S U23051 ( .I(gray_img[765]), .O(n26340) );
  MOAI1S U23052 ( .A1(n16003), .A2(n26340), .B1(n15866), .B2(gray_img[2029]), 
        .O(n17138) );
  AN4B1S U23053 ( .I1(n17141), .I2(n17140), .I3(n17139), .B1(n17138), .O(
        n17147) );
  AOI22S U23054 ( .A1(n15876), .A2(gray_img[1781]), .B1(n16188), .B2(
        gray_img[1277]), .O(n17146) );
  AOI22S U23055 ( .A1(n17778), .A2(gray_img[493]), .B1(n15895), .B2(
        gray_img[1533]), .O(n17145) );
  AOI22S U23056 ( .A1(n17591), .A2(gray_img[381]), .B1(gray_img[109]), .B2(
        n17779), .O(n17143) );
  AOI22S U23057 ( .A1(n15877), .A2(gray_img[365]), .B1(n15899), .B2(
        gray_img[749]), .O(n17142) );
  ND2S U23058 ( .I1(n17143), .I2(n17142), .O(n17144) );
  AN4B1S U23059 ( .I1(n17147), .I2(n17146), .I3(n17145), .B1(n17144), .O(
        n17160) );
  AOI22S U23060 ( .A1(n15874), .A2(gray_img[1133]), .B1(n17148), .B2(
        gray_img[1405]), .O(n17152) );
  AOI22S U23061 ( .A1(n16001), .A2(gray_img[757]), .B1(n15875), .B2(
        gray_img[125]), .O(n17151) );
  AOI22S U23062 ( .A1(n17807), .A2(gray_img[1013]), .B1(n15951), .B2(
        gray_img[1269]), .O(n17150) );
  INV1S U23063 ( .I(gray_img[253]), .O(n27564) );
  MOAI1S U23064 ( .A1(n17533), .A2(n27564), .B1(n17805), .B2(gray_img[1773]), 
        .O(n17149) );
  AN4B1S U23065 ( .I1(n17152), .I2(n17151), .I3(n17150), .B1(n17149), .O(
        n17158) );
  AOI22S U23066 ( .A1(n17795), .A2(gray_img[1005]), .B1(n17796), .B2(
        gray_img[1389]), .O(n17157) );
  AOI22S U23067 ( .A1(n15897), .A2(gray_img[2037]), .B1(n17797), .B2(
        gray_img[1517]), .O(n17156) );
  AOI22S U23068 ( .A1(n17605), .A2(gray_img[1141]), .B1(n15879), .B2(
        gray_img[1021]), .O(n17154) );
  AOI22S U23069 ( .A1(n17798), .A2(gray_img[373]), .B1(n15950), .B2(
        gray_img[245]), .O(n17153) );
  ND2S U23070 ( .I1(n17154), .I2(n17153), .O(n17155) );
  AN4B1S U23071 ( .I1(n17158), .I2(n17157), .I3(n17156), .B1(n17155), .O(
        n17159) );
  ND3S U23072 ( .I1(n17161), .I2(n17160), .I3(n17159), .O(n17162) );
  AOI22S U23073 ( .A1(n17163), .A2(n17817), .B1(n17819), .B2(n17162), .O(
        n17164) );
  ND2S U23074 ( .I1(n17165), .I2(n17164), .O(n17166) );
  NR2 U23075 ( .I1(n15995), .I2(n17957), .O(n17167) );
  NR2 U23076 ( .I1(n15994), .I2(n17973), .O(n17959) );
  NR2 U23077 ( .I1(n15995), .I2(n15871), .O(n17958) );
  NR2 U23078 ( .I1(n15996), .I2(n17957), .O(n17956) );
  NR2 U23079 ( .I1(n15997), .I2(n15943), .O(n17955) );
  FA1 U23080 ( .A(cro_mac[10]), .B(n17171), .CI(n17170), .CO(n17954), .S(
        n17367) );
  AOI22S U23081 ( .A1(n15913), .A2(gray_img[1474]), .B1(n17750), .B2(
        gray_img[450]), .O(n17175) );
  AOI22S U23082 ( .A1(n16000), .A2(gray_img[1090]), .B1(n17751), .B2(
        gray_img[1602]), .O(n17174) );
  AOI22S U23083 ( .A1(n15909), .A2(gray_img[194]), .B1(n15903), .B2(
        gray_img[1346]), .O(n17173) );
  INV1S U23084 ( .I(gray_img[1986]), .O(n23550) );
  MOAI1S U23085 ( .A1(n17753), .A2(n23550), .B1(n17752), .B2(gray_img[322]), 
        .O(n17172) );
  AN4B1S U23086 ( .I1(n17175), .I2(n17174), .I3(n17173), .B1(n17172), .O(
        n17192) );
  AOI22S U23087 ( .A1(n15902), .A2(gray_img[1730]), .B1(n17478), .B2(
        gray_img[66]), .O(n17179) );
  AOI22S U23088 ( .A1(n17758), .A2(gray_img[834]), .B1(n16165), .B2(
        gray_img[578]), .O(n17178) );
  AOI22S U23089 ( .A1(n17759), .A2(gray_img[1218]), .B1(n15901), .B2(
        gray_img[1858]), .O(n17177) );
  INV1S U23090 ( .I(gray_img[706]), .O(n27136) );
  MOAI1S U23091 ( .A1(n17760), .A2(n27136), .B1(n15900), .B2(gray_img[962]), 
        .O(n17176) );
  AN4B1S U23092 ( .I1(n17179), .I2(n17178), .I3(n17177), .B1(n17176), .O(
        n17191) );
  AOI22S U23093 ( .A1(n16116), .A2(gray_img[474]), .B1(n15914), .B2(
        gray_img[1754]), .O(n17183) );
  AOI22S U23094 ( .A1(n17770), .A2(gray_img[466]), .B1(n15873), .B2(
        gray_img[2010]), .O(n17182) );
  AOI22S U23095 ( .A1(n15917), .A2(gray_img[850]), .B1(n17765), .B2(
        gray_img[1866]), .O(n17181) );
  INV1S U23096 ( .I(gray_img[1618]), .O(n25514) );
  MOAI1S U23097 ( .A1(n17704), .A2(n25514), .B1(n17703), .B2(gray_img[602]), 
        .O(n17180) );
  AN4B1S U23098 ( .I1(n17183), .I2(n17182), .I3(n17181), .B1(n17180), .O(
        n17190) );
  INV1S U23099 ( .I(gray_img[594]), .O(n27015) );
  MOAI1S U23100 ( .A1(n17505), .A2(n27015), .B1(n16137), .B2(gray_img[842]), 
        .O(n17185) );
  INV1S U23101 ( .I(gray_img[1610]), .O(n25656) );
  MOAI1S U23102 ( .A1(n17381), .A2(n25656), .B1(n15908), .B2(gray_img[1626]), 
        .O(n17184) );
  NR2 U23103 ( .I1(n17185), .I2(n17184), .O(n17188) );
  AOI22S U23104 ( .A1(n15898), .A2(gray_img[858]), .B1(n15911), .B2(
        gray_img[1882]), .O(n17187) );
  AOI22S U23105 ( .A1(n15948), .A2(gray_img[1874]), .B1(n17709), .B2(
        gray_img[586]), .O(n17186) );
  ND3S U23106 ( .I1(n17188), .I2(n17187), .I3(n17186), .O(n17189) );
  AN4B1S U23107 ( .I1(n17192), .I2(n17191), .I3(n17190), .B1(n17189), .O(
        n17216) );
  AOI22S U23108 ( .A1(n15872), .A2(gray_img[1114]), .B1(n17785), .B2(
        gray_img[1226]), .O(n17196) );
  AOI22S U23109 ( .A1(n15878), .A2(gray_img[1362]), .B1(n17787), .B2(
        gray_img[202]), .O(n17195) );
  AOI22S U23110 ( .A1(n17329), .A2(gray_img[82]), .B1(n15949), .B2(
        gray_img[1490]), .O(n17194) );
  INV1S U23111 ( .I(gray_img[1994]), .O(n23563) );
  MOAI1S U23112 ( .A1(n15894), .A2(n23563), .B1(n17786), .B2(gray_img[730]), 
        .O(n17193) );
  AN4B1S U23113 ( .I1(n17196), .I2(n17195), .I3(n17194), .B1(n17193), .O(
        n17203) );
  AOI22S U23114 ( .A1(n15876), .A2(gray_img[1746]), .B1(n16188), .B2(
        gray_img[1242]), .O(n17202) );
  AOI22S U23115 ( .A1(n17778), .A2(gray_img[458]), .B1(n15895), .B2(
        gray_img[1498]), .O(n17201) );
  AOI22S U23116 ( .A1(n17197), .A2(gray_img[346]), .B1(n17779), .B2(
        gray_img[74]), .O(n17199) );
  AOI22S U23117 ( .A1(n15877), .A2(gray_img[330]), .B1(n15899), .B2(
        gray_img[714]), .O(n17198) );
  ND2S U23118 ( .I1(n17199), .I2(n17198), .O(n17200) );
  AN4B1S U23119 ( .I1(n17203), .I2(n17202), .I3(n17201), .B1(n17200), .O(
        n17215) );
  AOI22S U23120 ( .A1(n15897), .A2(gray_img[2002]), .B1(n17797), .B2(
        gray_img[1482]), .O(n17207) );
  AOI22S U23121 ( .A1(n17605), .A2(gray_img[1106]), .B1(n15879), .B2(
        gray_img[986]), .O(n17206) );
  AOI22S U23122 ( .A1(n17606), .A2(gray_img[338]), .B1(n15950), .B2(
        gray_img[210]), .O(n17205) );
  INV1S U23123 ( .I(gray_img[970]), .O(n22973) );
  MOAI1S U23124 ( .A1(n17718), .A2(n22973), .B1(n17796), .B2(gray_img[1354]), 
        .O(n17204) );
  AN4B1S U23125 ( .I1(n17207), .I2(n17206), .I3(n17205), .B1(n17204), .O(
        n17213) );
  AOI22S U23126 ( .A1(n16001), .A2(gray_img[722]), .B1(n15875), .B2(
        gray_img[90]), .O(n17212) );
  AOI22S U23127 ( .A1(n17723), .A2(gray_img[1098]), .B1(n17804), .B2(
        gray_img[1370]), .O(n17211) );
  AOI22S U23128 ( .A1(n17806), .A2(gray_img[218]), .B1(n17805), .B2(
        gray_img[1738]), .O(n17209) );
  AOI22S U23129 ( .A1(n17807), .A2(gray_img[978]), .B1(n15951), .B2(
        gray_img[1234]), .O(n17208) );
  ND2S U23130 ( .I1(n17209), .I2(n17208), .O(n17210) );
  AN4B1S U23131 ( .I1(n17213), .I2(n17212), .I3(n17211), .B1(n17210), .O(
        n17214) );
  ND3S U23132 ( .I1(n17216), .I2(n17215), .I3(n17214), .O(n17263) );
  AOI22S U23133 ( .A1(n15908), .A2(gray_img[1562]), .B1(n17743), .B2(
        gray_img[1546]), .O(n17220) );
  AOI22S U23134 ( .A1(n15898), .A2(gray_img[794]), .B1(n15911), .B2(
        gray_img[1818]), .O(n17219) );
  AOI22S U23135 ( .A1(n15948), .A2(gray_img[1810]), .B1(n17709), .B2(
        gray_img[522]), .O(n17218) );
  MOAI1S U23136 ( .A1(n17505), .A2(intadd_132_B_1_), .B1(n16137), .B2(
        gray_img[778]), .O(n17217) );
  AN4B1S U23137 ( .I1(n17220), .I2(n17219), .I3(n17218), .B1(n17217), .O(
        n17238) );
  AOI22S U23138 ( .A1(n16116), .A2(gray_img[410]), .B1(n15914), .B2(
        gray_img[1690]), .O(n17225) );
  AOI22S U23139 ( .A1(n17703), .A2(gray_img[538]), .B1(n17767), .B2(
        gray_img[1554]), .O(n17224) );
  AOI22S U23140 ( .A1(n15917), .A2(gray_img[786]), .B1(n17765), .B2(
        gray_img[1802]), .O(n17223) );
  INV1S U23141 ( .I(gray_img[402]), .O(n28736) );
  MOAI1S U23142 ( .A1(n17221), .A2(n28736), .B1(n15873), .B2(gray_img[1946]), 
        .O(n17222) );
  AN4B1S U23143 ( .I1(n17225), .I2(n17224), .I3(n17223), .B1(n17222), .O(
        n17237) );
  AOI22S U23144 ( .A1(n17752), .A2(gray_img[258]), .B1(n17696), .B2(
        gray_img[1922]), .O(n17229) );
  AOI22S U23145 ( .A1(n15913), .A2(gray_img[1410]), .B1(n17750), .B2(
        gray_img[386]), .O(n17228) );
  AOI22S U23146 ( .A1(n15909), .A2(gray_img[130]), .B1(n15903), .B2(
        gray_img[1282]), .O(n17227) );
  INV1S U23147 ( .I(gray_img[1538]), .O(n26590) );
  MOAI1S U23148 ( .A1(n15942), .A2(n26590), .B1(n16000), .B2(gray_img[1026]), 
        .O(n17226) );
  AN4B1S U23149 ( .I1(n17229), .I2(n17228), .I3(n17227), .B1(n17226), .O(
        n17236) );
  INV1S U23150 ( .I(gray_img[514]), .O(n29919) );
  MOAI1S U23151 ( .A1(n17640), .A2(n29919), .B1(n17758), .B2(gray_img[770]), 
        .O(n17231) );
  INV1S U23152 ( .I(gray_img[1154]), .O(n26629) );
  MOAI1S U23153 ( .A1(n17518), .A2(n26629), .B1(n15901), .B2(gray_img[1794]), 
        .O(n17230) );
  NR2 U23154 ( .I1(n17231), .I2(n17230), .O(n17234) );
  AOI22S U23155 ( .A1(n15900), .A2(gray_img[898]), .B1(n17639), .B2(
        gray_img[642]), .O(n17233) );
  AOI22S U23156 ( .A1(n15902), .A2(gray_img[1666]), .B1(n15912), .B2(
        gray_img[2]), .O(n17232) );
  ND3S U23157 ( .I1(n17234), .I2(n17233), .I3(n17232), .O(n17235) );
  AN4B1S U23158 ( .I1(n17238), .I2(n17237), .I3(n17236), .B1(n17235), .O(
        n17261) );
  AOI22S U23159 ( .A1(n15872), .A2(gray_img[1050]), .B1(n17785), .B2(
        gray_img[1162]), .O(n17242) );
  AOI22S U23160 ( .A1(n15878), .A2(gray_img[1298]), .B1(n17787), .B2(
        gray_img[138]), .O(n17241) );
  AOI22S U23161 ( .A1(n17329), .A2(gray_img[18]), .B1(n15949), .B2(
        gray_img[1426]), .O(n17240) );
  INV1S U23162 ( .I(gray_img[1930]), .O(n29402) );
  MOAI1S U23163 ( .A1(n15894), .A2(n29402), .B1(n17786), .B2(gray_img[666]), 
        .O(n17239) );
  AN4B1S U23164 ( .I1(n17242), .I2(n17241), .I3(n17240), .B1(n17239), .O(
        n17248) );
  AOI22S U23165 ( .A1(n15876), .A2(gray_img[1682]), .B1(n16188), .B2(
        gray_img[1178]), .O(n17247) );
  AOI22S U23166 ( .A1(n17778), .A2(gray_img[394]), .B1(n15895), .B2(
        gray_img[1434]), .O(n17246) );
  AOI22S U23167 ( .A1(n17591), .A2(gray_img[282]), .B1(n17779), .B2(
        gray_img[10]), .O(n17244) );
  AOI22S U23168 ( .A1(n15877), .A2(gray_img[266]), .B1(n16368), .B2(
        gray_img[650]), .O(n17243) );
  ND2S U23169 ( .I1(n17244), .I2(n17243), .O(n17245) );
  AN4B1S U23170 ( .I1(n17248), .I2(n17247), .I3(n17246), .B1(n17245), .O(
        n17260) );
  AOI22S U23171 ( .A1(n15897), .A2(gray_img[1938]), .B1(n17797), .B2(
        gray_img[1418]), .O(n17252) );
  AOI22S U23172 ( .A1(n17605), .A2(gray_img[1042]), .B1(n15879), .B2(
        gray_img[922]), .O(n17251) );
  AOI22S U23173 ( .A1(n17717), .A2(gray_img[274]), .B1(n15950), .B2(
        gray_img[146]), .O(n17250) );
  INV1S U23174 ( .I(gray_img[906]), .O(n29606) );
  MOAI1S U23175 ( .A1(n17718), .A2(n29606), .B1(n17796), .B2(gray_img[1290]), 
        .O(n17249) );
  AN4B1S U23176 ( .I1(n17252), .I2(n17251), .I3(n17250), .B1(n17249), .O(
        n17258) );
  AOI22S U23177 ( .A1(n16001), .A2(gray_img[658]), .B1(n15896), .B2(
        gray_img[26]), .O(n17257) );
  AOI22S U23178 ( .A1(n17723), .A2(gray_img[1034]), .B1(n17804), .B2(
        gray_img[1306]), .O(n17256) );
  AOI22S U23179 ( .A1(n17806), .A2(gray_img[154]), .B1(n17805), .B2(
        gray_img[1674]), .O(n17254) );
  AOI22S U23180 ( .A1(n17807), .A2(gray_img[914]), .B1(n15951), .B2(
        gray_img[1170]), .O(n17253) );
  ND2S U23181 ( .I1(n17254), .I2(n17253), .O(n17255) );
  AN4B1S U23182 ( .I1(n17258), .I2(n17257), .I3(n17256), .B1(n17255), .O(
        n17259) );
  ND3S U23183 ( .I1(n17261), .I2(n17260), .I3(n17259), .O(n17262) );
  AOI22S U23184 ( .A1(n17263), .A2(n17690), .B1(n17262), .B2(n17688), .O(
        n17356) );
  AOI22S U23185 ( .A1(n16116), .A2(gray_img[506]), .B1(n15914), .B2(
        gray_img[1786]), .O(n17267) );
  AOI22S U23186 ( .A1(n17703), .A2(gray_img[634]), .B1(n17767), .B2(
        gray_img[1650]), .O(n17266) );
  AOI22S U23187 ( .A1(n17770), .A2(gray_img[498]), .B1(n15873), .B2(
        gray_img[2042]), .O(n17265) );
  INV1S U23188 ( .I(gray_img[882]), .O(n26377) );
  MOAI1S U23189 ( .A1(n17766), .A2(n26377), .B1(n17765), .B2(gray_img[1898]), 
        .O(n17264) );
  AN4B1S U23190 ( .I1(n17267), .I2(n17266), .I3(n17265), .B1(n17264), .O(
        n17284) );
  AOI22S U23191 ( .A1(n15913), .A2(gray_img[1506]), .B1(n17750), .B2(
        gray_img[482]), .O(n17271) );
  AOI22S U23192 ( .A1(n16000), .A2(gray_img[1122]), .B1(n17751), .B2(
        gray_img[1634]), .O(n17270) );
  AOI22S U23193 ( .A1(n15909), .A2(gray_img[226]), .B1(n15903), .B2(
        gray_img[1378]), .O(n17269) );
  INV1S U23194 ( .I(gray_img[2018]), .O(n25838) );
  MOAI1S U23195 ( .A1(n17753), .A2(n25838), .B1(n17752), .B2(gray_img[354]), 
        .O(n17268) );
  AN4B1S U23196 ( .I1(n17271), .I2(n17270), .I3(n17269), .B1(n17268), .O(
        n17283) );
  AOI22S U23197 ( .A1(n15902), .A2(gray_img[1762]), .B1(n15912), .B2(
        gray_img[98]), .O(n17275) );
  AOI22S U23198 ( .A1(n17758), .A2(gray_img[866]), .B1(n16165), .B2(
        gray_img[610]), .O(n17274) );
  AOI22S U23199 ( .A1(n17759), .A2(gray_img[1250]), .B1(n15901), .B2(
        gray_img[1890]), .O(n17273) );
  INV1S U23200 ( .I(gray_img[738]), .O(n26164) );
  MOAI1S U23201 ( .A1(n17760), .A2(n26164), .B1(n15900), .B2(gray_img[994]), 
        .O(n17272) );
  AN4B1S U23202 ( .I1(n17275), .I2(n17274), .I3(n17273), .B1(n17272), .O(
        n17282) );
  INV1S U23203 ( .I(gray_img[890]), .O(n26390) );
  MOAI1S U23204 ( .A1(n15946), .A2(n26390), .B1(n15911), .B2(gray_img[1914]), 
        .O(n17277) );
  INV1S U23205 ( .I(gray_img[618]), .O(n26189) );
  MOAI1S U23206 ( .A1(n17745), .A2(n26189), .B1(n15948), .B2(gray_img[1906]), 
        .O(n17276) );
  NR2 U23207 ( .I1(n17277), .I2(n17276), .O(n17280) );
  AOI22S U23208 ( .A1(n15908), .A2(gray_img[1658]), .B1(n17743), .B2(
        gray_img[1642]), .O(n17279) );
  AOI22S U23209 ( .A1(n16137), .A2(gray_img[874]), .B1(n17744), .B2(
        gray_img[626]), .O(n17278) );
  ND3S U23210 ( .I1(n17280), .I2(n17279), .I3(n17278), .O(n17281) );
  AOI22S U23211 ( .A1(n15872), .A2(gray_img[1146]), .B1(n17785), .B2(
        gray_img[1258]), .O(n17288) );
  AOI22S U23212 ( .A1(n15878), .A2(gray_img[1394]), .B1(n17787), .B2(
        gray_img[234]), .O(n17287) );
  AOI22S U23213 ( .A1(n17329), .A2(gray_img[114]), .B1(n15949), .B2(
        gray_img[1522]), .O(n17286) );
  INV1S U23214 ( .I(gray_img[2026]), .O(n25850) );
  MOAI1S U23215 ( .A1(n15894), .A2(n25850), .B1(n17786), .B2(gray_img[762]), 
        .O(n17285) );
  AN4B1S U23216 ( .I1(n17288), .I2(n17287), .I3(n17286), .B1(n17285), .O(
        n17294) );
  AOI22S U23217 ( .A1(n15876), .A2(gray_img[1778]), .B1(n16188), .B2(
        gray_img[1274]), .O(n17293) );
  AOI22S U23218 ( .A1(n17778), .A2(gray_img[490]), .B1(n15895), .B2(
        gray_img[1530]), .O(n17292) );
  AOI22S U23219 ( .A1(n17591), .A2(gray_img[378]), .B1(n17779), .B2(
        gray_img[106]), .O(n17290) );
  AOI22S U23220 ( .A1(n15877), .A2(gray_img[362]), .B1(n15899), .B2(
        gray_img[746]), .O(n17289) );
  ND2S U23221 ( .I1(n17290), .I2(n17289), .O(n17291) );
  AN4B1S U23222 ( .I1(n17294), .I2(n17293), .I3(n17292), .B1(n17291), .O(
        n17306) );
  AOI22S U23223 ( .A1(n15874), .A2(gray_img[1130]), .B1(n17804), .B2(
        gray_img[1402]), .O(n17298) );
  AOI22S U23224 ( .A1(n16001), .A2(gray_img[754]), .B1(n15875), .B2(
        gray_img[122]), .O(n17297) );
  AOI22S U23225 ( .A1(n17807), .A2(gray_img[1010]), .B1(n15951), .B2(
        gray_img[1266]), .O(n17296) );
  INV1S U23226 ( .I(gray_img[250]), .O(n27558) );
  MOAI1S U23227 ( .A1(n17533), .A2(n27558), .B1(n17805), .B2(gray_img[1770]), 
        .O(n17295) );
  AN4B1S U23228 ( .I1(n17298), .I2(n17297), .I3(n17296), .B1(n17295), .O(
        n17304) );
  AOI22S U23229 ( .A1(n17796), .A2(gray_img[1386]), .B1(n17795), .B2(
        gray_img[1002]), .O(n17303) );
  AOI22S U23230 ( .A1(n17716), .A2(gray_img[2034]), .B1(n17797), .B2(
        gray_img[1514]), .O(n17302) );
  AOI22S U23231 ( .A1(n17605), .A2(gray_img[1138]), .B1(n15879), .B2(
        gray_img[1018]), .O(n17300) );
  AOI22S U23232 ( .A1(n17606), .A2(gray_img[370]), .B1(n15950), .B2(
        gray_img[242]), .O(n17299) );
  ND2S U23233 ( .I1(n17300), .I2(n17299), .O(n17301) );
  AN4B1S U23234 ( .I1(n17304), .I2(n17303), .I3(n17302), .B1(n17301), .O(
        n17305) );
  ND3S U23235 ( .I1(n17307), .I2(n17306), .I3(n17305), .O(n17354) );
  AOI22S U23236 ( .A1(n15908), .A2(gray_img[1594]), .B1(n17743), .B2(
        gray_img[1578]), .O(n17311) );
  AOI22S U23237 ( .A1(n15898), .A2(gray_img[826]), .B1(n15911), .B2(
        gray_img[1850]), .O(n17310) );
  AOI22S U23238 ( .A1(n16137), .A2(gray_img[810]), .B1(n17744), .B2(
        gray_img[562]), .O(n17309) );
  INV1S U23239 ( .I(gray_img[554]), .O(n28609) );
  MOAI1S U23240 ( .A1(n17745), .A2(n28609), .B1(n15948), .B2(gray_img[1842]), 
        .O(n17308) );
  AN4B1S U23241 ( .I1(n17311), .I2(n17310), .I3(n17309), .B1(n17308), .O(
        n17328) );
  AOI22S U23242 ( .A1(n16116), .A2(gray_img[442]), .B1(n15914), .B2(
        gray_img[1722]), .O(n17315) );
  AOI22S U23243 ( .A1(n17703), .A2(gray_img[570]), .B1(n17767), .B2(
        gray_img[1586]), .O(n17314) );
  AOI22S U23244 ( .A1(n17770), .A2(gray_img[434]), .B1(n15873), .B2(
        gray_img[1978]), .O(n17313) );
  INV1S U23245 ( .I(gray_img[818]), .O(n26100) );
  MOAI1S U23246 ( .A1(n17766), .A2(n26100), .B1(n17765), .B2(gray_img[1834]), 
        .O(n17312) );
  AN4B1S U23247 ( .I1(n17315), .I2(n17314), .I3(n17313), .B1(n17312), .O(
        n17327) );
  AOI22S U23248 ( .A1(n15913), .A2(gray_img[1442]), .B1(n17750), .B2(
        gray_img[418]), .O(n17319) );
  AOI22S U23249 ( .A1(n16000), .A2(gray_img[1058]), .B1(n17751), .B2(
        gray_img[1570]), .O(n17318) );
  AOI22S U23250 ( .A1(n15909), .A2(gray_img[162]), .B1(n15903), .B2(
        gray_img[1314]), .O(n17317) );
  INV1S U23251 ( .I(gray_img[1954]), .O(n26658) );
  MOAI1S U23252 ( .A1(n17753), .A2(n26658), .B1(n17752), .B2(gray_img[290]), 
        .O(n17316) );
  AN4B1S U23253 ( .I1(n17319), .I2(n17318), .I3(n17317), .B1(n17316), .O(
        n17326) );
  INV1S U23254 ( .I(gray_img[546]), .O(n28622) );
  MOAI1S U23255 ( .A1(n17640), .A2(n28622), .B1(n17758), .B2(gray_img[802]), 
        .O(n17321) );
  INV1S U23256 ( .I(gray_img[1186]), .O(n23010) );
  MOAI1S U23257 ( .A1(n17518), .A2(n23010), .B1(n15901), .B2(gray_img[1826]), 
        .O(n17320) );
  NR2 U23258 ( .I1(n17321), .I2(n17320), .O(n17324) );
  AOI22S U23259 ( .A1(n15900), .A2(gray_img[930]), .B1(n17639), .B2(
        gray_img[674]), .O(n17323) );
  AOI22S U23260 ( .A1(n15902), .A2(gray_img[1698]), .B1(n17478), .B2(
        gray_img[34]), .O(n17322) );
  ND3S U23261 ( .I1(n17324), .I2(n17323), .I3(n17322), .O(n17325) );
  AN4B1S U23262 ( .I1(n17328), .I2(n17327), .I3(n17326), .B1(n17325), .O(
        n17352) );
  AOI22S U23263 ( .A1(n15872), .A2(gray_img[1082]), .B1(n17785), .B2(
        gray_img[1194]), .O(n17333) );
  AOI22S U23264 ( .A1(n15878), .A2(gray_img[1330]), .B1(n17787), .B2(
        gray_img[170]), .O(n17332) );
  AOI22S U23265 ( .A1(n17329), .A2(gray_img[50]), .B1(n15949), .B2(
        gray_img[1458]), .O(n17331) );
  INV1S U23266 ( .I(gray_img[1962]), .O(n26671) );
  MOAI1S U23267 ( .A1(n15894), .A2(n26671), .B1(n17786), .B2(gray_img[698]), 
        .O(n17330) );
  AN4B1S U23268 ( .I1(n17333), .I2(n17332), .I3(n17331), .B1(n17330), .O(
        n17339) );
  AOI22S U23269 ( .A1(n15876), .A2(gray_img[1714]), .B1(n16188), .B2(
        gray_img[1210]), .O(n17338) );
  AOI22S U23270 ( .A1(n17778), .A2(gray_img[426]), .B1(n15895), .B2(
        gray_img[1466]), .O(n17337) );
  AOI22S U23271 ( .A1(n17780), .A2(gray_img[314]), .B1(n17779), .B2(
        gray_img[42]), .O(n17335) );
  AOI22S U23272 ( .A1(n15877), .A2(gray_img[298]), .B1(n16368), .B2(
        gray_img[682]), .O(n17334) );
  ND2S U23273 ( .I1(n17335), .I2(n17334), .O(n17336) );
  AN4B1S U23274 ( .I1(n17339), .I2(n17338), .I3(n17337), .B1(n17336), .O(
        n17351) );
  AOI22S U23275 ( .A1(n15897), .A2(gray_img[1970]), .B1(n17797), .B2(
        gray_img[1450]), .O(n17343) );
  AOI22S U23276 ( .A1(n17605), .A2(gray_img[1074]), .B1(n15879), .B2(
        gray_img[954]), .O(n17342) );
  AOI22S U23277 ( .A1(n17606), .A2(gray_img[306]), .B1(n15950), .B2(
        gray_img[178]), .O(n17341) );
  INV1S U23278 ( .I(gray_img[938]), .O(n23210) );
  MOAI1S U23279 ( .A1(n17718), .A2(n23210), .B1(n17796), .B2(gray_img[1322]), 
        .O(n17340) );
  AN4B1S U23280 ( .I1(n17343), .I2(n17342), .I3(n17341), .B1(n17340), .O(
        n17349) );
  AOI22S U23281 ( .A1(n16001), .A2(gray_img[690]), .B1(n15875), .B2(
        gray_img[58]), .O(n17348) );
  AOI22S U23282 ( .A1(n17723), .A2(gray_img[1066]), .B1(n17804), .B2(
        gray_img[1338]), .O(n17347) );
  AOI22S U23283 ( .A1(n17806), .A2(gray_img[186]), .B1(n17805), .B2(
        gray_img[1706]), .O(n17345) );
  AOI22S U23284 ( .A1(n17807), .A2(gray_img[946]), .B1(n15951), .B2(
        gray_img[1202]), .O(n17344) );
  ND2S U23285 ( .I1(n17345), .I2(n17344), .O(n17346) );
  AN4B1S U23286 ( .I1(n17349), .I2(n17348), .I3(n17347), .B1(n17346), .O(
        n17350) );
  ND3S U23287 ( .I1(n17352), .I2(n17351), .I3(n17350), .O(n17353) );
  AOI22S U23288 ( .A1(n17354), .A2(n17819), .B1(n17353), .B2(n17817), .O(
        n17355) );
  ND2S U23289 ( .I1(n17356), .I2(n17355), .O(n17357) );
  INV2 U23290 ( .I(n17357), .O(n17868) );
  NR2 U23291 ( .I1(n15997), .I2(n17868), .O(n17559) );
  NR2 U23292 ( .I1(n15994), .I2(n17957), .O(n17558) );
  AO222S U23293 ( .A1(template_reg[9]), .A2(n17581), .B1(template_reg[1]), 
        .B2(n17579), .C1(n17580), .C2(template_reg[17]), .O(n17363) );
  ND2S U23294 ( .I1(n17358), .I2(cnt_cro_3b3[0]), .O(n17361) );
  AOI22S U23295 ( .A1(n17584), .A2(template_reg[65]), .B1(n17583), .B2(
        template_reg[57]), .O(n17360) );
  ND2S U23296 ( .I1(n17585), .I2(template_reg[49]), .O(n17359) );
  NR2 U23297 ( .I1(n15991), .I2(n17973), .O(n17563) );
  NR2 U23298 ( .I1(n15995), .I2(n15943), .O(n17562) );
  NR2 U23299 ( .I1(n15996), .I2(n17873), .O(n17561) );
  FA1 U23300 ( .A(cro_mac[9]), .B(n17365), .CI(n17364), .CO(n17368), .S(n17560) );
  FA1 U23301 ( .A(n17368), .B(n17367), .CI(n17366), .CO(n17965), .S(n17570) );
  NR2 U23302 ( .I1(n15995), .I2(n17873), .O(n17847) );
  NR2 U23303 ( .I1(n15993), .I2(n17957), .O(n17846) );
  AOI22S U23304 ( .A1(n15913), .A2(gray_img[1473]), .B1(n17750), .B2(
        gray_img[449]), .O(n17372) );
  AOI22S U23305 ( .A1(n16000), .A2(gray_img[1089]), .B1(n17751), .B2(
        gray_img[1601]), .O(n17371) );
  AOI22S U23306 ( .A1(n15909), .A2(gray_img[193]), .B1(n15903), .B2(
        gray_img[1345]), .O(n17370) );
  MOAI1S U23307 ( .A1(n17753), .A2(intadd_25_B_0_), .B1(n17752), .B2(
        gray_img[321]), .O(n17369) );
  AN4B1S U23308 ( .I1(n17372), .I2(n17371), .I3(n17370), .B1(n17369), .O(
        n17390) );
  AOI22S U23309 ( .A1(n15902), .A2(gray_img[1729]), .B1(n17478), .B2(
        gray_img[65]), .O(n17376) );
  AOI22S U23310 ( .A1(n17758), .A2(gray_img[833]), .B1(n16165), .B2(
        gray_img[577]), .O(n17375) );
  AOI22S U23311 ( .A1(n17759), .A2(gray_img[1217]), .B1(n15901), .B2(
        gray_img[1857]), .O(n17374) );
  MOAI1S U23312 ( .A1(n17760), .A2(intadd_109_CI), .B1(n15900), .B2(
        gray_img[961]), .O(n17373) );
  AN4B1S U23313 ( .I1(n17376), .I2(n17375), .I3(n17374), .B1(n17373), .O(
        n17389) );
  AOI22S U23314 ( .A1(n16116), .A2(gray_img[473]), .B1(n15914), .B2(
        gray_img[1753]), .O(n17380) );
  AOI22S U23315 ( .A1(n17770), .A2(gray_img[465]), .B1(n15873), .B2(
        gray_img[2009]), .O(n17379) );
  AOI22S U23316 ( .A1(n15917), .A2(gray_img[849]), .B1(n17765), .B2(
        gray_img[1865]), .O(n17378) );
  INV1S U23317 ( .I(gray_img[1617]), .O(n25512) );
  MOAI1S U23318 ( .A1(n17704), .A2(n25512), .B1(n17703), .B2(gray_img[601]), 
        .O(n17377) );
  AN4B1S U23319 ( .I1(n17380), .I2(n17379), .I3(n17378), .B1(n17377), .O(
        n17388) );
  MOAI1S U23320 ( .A1(n17505), .A2(intadd_105_CI), .B1(n16137), .B2(
        gray_img[841]), .O(n17383) );
  INV1S U23321 ( .I(gray_img[1609]), .O(n25654) );
  MOAI1S U23322 ( .A1(n17381), .A2(n25654), .B1(n15908), .B2(gray_img[1625]), 
        .O(n17382) );
  NR2 U23323 ( .I1(n17383), .I2(n17382), .O(n17386) );
  AOI22S U23324 ( .A1(n15898), .A2(gray_img[857]), .B1(n15911), .B2(
        gray_img[1881]), .O(n17385) );
  AOI22S U23325 ( .A1(n15948), .A2(gray_img[1873]), .B1(n17709), .B2(
        gray_img[585]), .O(n17384) );
  ND3S U23326 ( .I1(n17386), .I2(n17385), .I3(n17384), .O(n17387) );
  AN4B1S U23327 ( .I1(n17390), .I2(n17389), .I3(n17388), .B1(n17387), .O(
        n17413) );
  AOI22S U23328 ( .A1(n17778), .A2(gray_img[457]), .B1(n15895), .B2(
        gray_img[1497]), .O(n17394) );
  AOI22S U23329 ( .A1(n15877), .A2(gray_img[329]), .B1(n15899), .B2(
        gray_img[713]), .O(n17393) );
  AOI22S U23330 ( .A1(n15876), .A2(gray_img[1745]), .B1(n16188), .B2(
        gray_img[1241]), .O(n17392) );
  MOAI1S U23331 ( .A1(n16002), .A2(intadd_130_B_0_), .B1(n17780), .B2(
        gray_img[345]), .O(n17391) );
  AN4B1S U23332 ( .I1(n17394), .I2(n17393), .I3(n17392), .B1(n17391), .O(
        n17411) );
  AOI22S U23333 ( .A1(n15872), .A2(gray_img[1113]), .B1(n17785), .B2(
        gray_img[1225]), .O(n17398) );
  AOI22S U23334 ( .A1(n15878), .A2(gray_img[1361]), .B1(n17787), .B2(
        gray_img[201]), .O(n17397) );
  INV2 U23335 ( .I(n15941), .O(n17788) );
  AOI22S U23336 ( .A1(n17788), .A2(gray_img[81]), .B1(n15949), .B2(
        gray_img[1489]), .O(n17396) );
  INV1S U23337 ( .I(gray_img[1993]), .O(n23561) );
  MOAI1S U23338 ( .A1(n15894), .A2(n23561), .B1(n17786), .B2(gray_img[729]), 
        .O(n17395) );
  AN4B1S U23339 ( .I1(n17398), .I2(n17397), .I3(n17396), .B1(n17395), .O(
        n17410) );
  AOI22S U23340 ( .A1(n15897), .A2(gray_img[2001]), .B1(n17797), .B2(
        gray_img[1481]), .O(n17402) );
  AOI22S U23341 ( .A1(n17605), .A2(gray_img[1105]), .B1(n15879), .B2(
        gray_img[985]), .O(n17401) );
  AOI22S U23342 ( .A1(n17606), .A2(gray_img[337]), .B1(n15950), .B2(
        gray_img[209]), .O(n17400) );
  MOAI1S U23343 ( .A1(n17718), .A2(intadd_98_CI), .B1(n17796), .B2(
        gray_img[1353]), .O(n17399) );
  AN4B1S U23344 ( .I1(n17402), .I2(n17401), .I3(n17400), .B1(n17399), .O(
        n17409) );
  MOAI1S U23345 ( .A1(n15868), .A2(intadd_188_B_0_), .B1(n16001), .B2(
        gray_img[721]), .O(n17404) );
  INV1S U23346 ( .I(gray_img[1369]), .O(n28360) );
  MOAI1S U23347 ( .A1(n17660), .A2(n28360), .B1(n15874), .B2(gray_img[1097]), 
        .O(n17403) );
  NR2 U23348 ( .I1(n17404), .I2(n17403), .O(n17407) );
  AOI22S U23349 ( .A1(n17807), .A2(gray_img[977]), .B1(n15951), .B2(
        gray_img[1233]), .O(n17406) );
  AOI22S U23350 ( .A1(n17806), .A2(gray_img[217]), .B1(n17805), .B2(
        gray_img[1737]), .O(n17405) );
  ND3S U23351 ( .I1(n17407), .I2(n17406), .I3(n17405), .O(n17408) );
  AN4B1S U23352 ( .I1(n17411), .I2(n17410), .I3(n17409), .B1(n17408), .O(
        n17412) );
  ND2S U23353 ( .I1(n17413), .I2(n17412), .O(n17459) );
  AOI22S U23354 ( .A1(n15908), .A2(gray_img[1593]), .B1(n17743), .B2(
        gray_img[1577]), .O(n17417) );
  AOI22S U23355 ( .A1(n15898), .A2(gray_img[825]), .B1(n15911), .B2(
        gray_img[1849]), .O(n17416) );
  AOI22S U23356 ( .A1(n16137), .A2(gray_img[809]), .B1(n17744), .B2(
        gray_img[561]), .O(n17415) );
  MOAI1S U23357 ( .A1(n17745), .A2(intadd_137_B_0_), .B1(n15948), .B2(
        gray_img[1841]), .O(n17414) );
  AN4B1S U23358 ( .I1(n17417), .I2(n17416), .I3(n17415), .B1(n17414), .O(
        n17434) );
  AOI22S U23359 ( .A1(n16116), .A2(gray_img[441]), .B1(n15914), .B2(
        gray_img[1721]), .O(n17421) );
  AOI22S U23360 ( .A1(n17770), .A2(gray_img[433]), .B1(n15873), .B2(
        gray_img[1977]), .O(n17420) );
  AOI22S U23361 ( .A1(n15917), .A2(gray_img[817]), .B1(n17765), .B2(
        gray_img[1833]), .O(n17419) );
  MOAI1S U23362 ( .A1(n17674), .A2(intadd_189_A_0_), .B1(n17767), .B2(
        gray_img[1585]), .O(n17418) );
  AN4B1S U23363 ( .I1(n17421), .I2(n17420), .I3(n17419), .B1(n17418), .O(
        n17433) );
  AOI22S U23364 ( .A1(n15913), .A2(gray_img[1441]), .B1(n17750), .B2(
        gray_img[417]), .O(n17425) );
  AOI22S U23365 ( .A1(n16000), .A2(gray_img[1057]), .B1(n17751), .B2(
        gray_img[1569]), .O(n17424) );
  AOI22S U23366 ( .A1(n15909), .A2(gray_img[161]), .B1(n15903), .B2(
        gray_img[1313]), .O(n17423) );
  INV1S U23367 ( .I(gray_img[1953]), .O(n26656) );
  MOAI1S U23368 ( .A1(n17753), .A2(n26656), .B1(n17752), .B2(gray_img[289]), 
        .O(n17422) );
  AN4B1S U23369 ( .I1(n17425), .I2(n17424), .I3(n17423), .B1(n17422), .O(
        n17432) );
  INV1S U23370 ( .I(gray_img[545]), .O(n28620) );
  MOAI1S U23371 ( .A1(n17640), .A2(n28620), .B1(n17758), .B2(gray_img[801]), 
        .O(n17427) );
  MOAI1S U23372 ( .A1(n17518), .A2(intadd_83_CI), .B1(n15901), .B2(
        gray_img[1825]), .O(n17426) );
  NR2 U23373 ( .I1(n17427), .I2(n17426), .O(n17430) );
  AOI22S U23374 ( .A1(n15900), .A2(gray_img[929]), .B1(n17639), .B2(
        gray_img[673]), .O(n17429) );
  AOI22S U23375 ( .A1(n15902), .A2(gray_img[1697]), .B1(n15912), .B2(
        gray_img[33]), .O(n17428) );
  ND3S U23376 ( .I1(n17430), .I2(n17429), .I3(n17428), .O(n17431) );
  AN4B1S U23377 ( .I1(n17434), .I2(n17433), .I3(n17432), .B1(n17431), .O(
        n17457) );
  AOI22S U23378 ( .A1(n15874), .A2(gray_img[1065]), .B1(n17804), .B2(
        gray_img[1337]), .O(n17438) );
  AOI22S U23379 ( .A1(n17806), .A2(gray_img[185]), .B1(n17805), .B2(
        gray_img[1705]), .O(n17437) );
  AOI22S U23380 ( .A1(n17807), .A2(gray_img[945]), .B1(n15951), .B2(
        gray_img[1201]), .O(n17436) );
  MOAI1S U23381 ( .A1(n15868), .A2(n27709), .B1(n16001), .B2(gray_img[689]), 
        .O(n17435) );
  AN4B1S U23382 ( .I1(n17438), .I2(n17437), .I3(n17436), .B1(n17435), .O(
        n17455) );
  AOI22S U23383 ( .A1(n15872), .A2(gray_img[1081]), .B1(n17785), .B2(
        gray_img[1193]), .O(n17442) );
  AOI22S U23384 ( .A1(n15878), .A2(gray_img[1329]), .B1(n17787), .B2(
        gray_img[169]), .O(n17441) );
  AOI22S U23385 ( .A1(n17788), .A2(gray_img[49]), .B1(n15949), .B2(
        gray_img[1457]), .O(n17440) );
  INV1S U23386 ( .I(gray_img[1961]), .O(n26669) );
  MOAI1S U23387 ( .A1(n15894), .A2(n26669), .B1(n17786), .B2(gray_img[697]), 
        .O(n17439) );
  AN4B1S U23388 ( .I1(n17442), .I2(n17441), .I3(n17440), .B1(n17439), .O(
        n17454) );
  AOI22S U23389 ( .A1(n15897), .A2(gray_img[1969]), .B1(n17797), .B2(
        gray_img[1449]), .O(n17446) );
  AOI22S U23390 ( .A1(n17605), .A2(gray_img[1073]), .B1(n15879), .B2(
        gray_img[953]), .O(n17445) );
  AOI22S U23391 ( .A1(n17717), .A2(gray_img[305]), .B1(n15950), .B2(
        gray_img[177]), .O(n17444) );
  MOAI1S U23392 ( .A1(n17718), .A2(intadd_162_CI), .B1(n17796), .B2(
        gray_img[1321]), .O(n17443) );
  AN4B1S U23393 ( .I1(n17446), .I2(n17445), .I3(n17444), .B1(n17443), .O(
        n17453) );
  MOAI1S U23394 ( .A1(n15947), .A2(intadd_44_CI), .B1(n16188), .B2(
        gray_img[1209]), .O(n17448) );
  MOAI1S U23395 ( .A1(n15867), .A2(intadd_134_CI), .B1(n17778), .B2(
        gray_img[425]), .O(n17447) );
  NR2 U23396 ( .I1(n17448), .I2(n17447), .O(n17451) );
  AOI22S U23397 ( .A1(n17780), .A2(gray_img[313]), .B1(n17779), .B2(
        gray_img[41]), .O(n17450) );
  AOI22S U23398 ( .A1(n15877), .A2(gray_img[297]), .B1(n15899), .B2(
        gray_img[681]), .O(n17449) );
  ND3S U23399 ( .I1(n17451), .I2(n17450), .I3(n17449), .O(n17452) );
  AN4B1S U23400 ( .I1(n17455), .I2(n17454), .I3(n17453), .B1(n17452), .O(
        n17456) );
  ND2S U23401 ( .I1(n17457), .I2(n17456), .O(n17458) );
  AOI22S U23402 ( .A1(n17459), .A2(n17690), .B1(n17458), .B2(n17817), .O(
        n17556) );
  AOI22S U23403 ( .A1(n15872), .A2(gray_img[1145]), .B1(n17785), .B2(
        gray_img[1257]), .O(n17463) );
  AOI22S U23404 ( .A1(n15878), .A2(gray_img[1393]), .B1(n17787), .B2(
        gray_img[233]), .O(n17462) );
  AOI22S U23405 ( .A1(n17788), .A2(gray_img[113]), .B1(n15949), .B2(
        gray_img[1521]), .O(n17461) );
  MOAI1S U23406 ( .A1(n15894), .A2(intadd_5_CI), .B1(n17786), .B2(
        gray_img[761]), .O(n17460) );
  AN4B1S U23407 ( .I1(n17463), .I2(n17462), .I3(n17461), .B1(n17460), .O(
        n17469) );
  INV1S U23408 ( .I(gray_img[1777]), .O(n25996) );
  MOAI1S U23409 ( .A1(n15947), .A2(n25996), .B1(n16188), .B2(gray_img[1273]), 
        .O(n17465) );
  MOAI1S U23410 ( .A1(n15867), .A2(intadd_145_CI), .B1(n17778), .B2(
        gray_img[489]), .O(n17464) );
  NR2 U23411 ( .I1(n17465), .I2(n17464), .O(n17468) );
  AOI22S U23412 ( .A1(n17591), .A2(gray_img[377]), .B1(n17779), .B2(
        gray_img[105]), .O(n17467) );
  INV1S U23413 ( .I(gray_img[361]), .O(n27451) );
  MOAI1S U23414 ( .A1(n16518), .A2(n27451), .B1(n15899), .B2(gray_img[745]), 
        .O(n17466) );
  AN4B1S U23415 ( .I1(n17469), .I2(n17468), .I3(n17467), .B1(n17466), .O(
        n17504) );
  AOI22S U23416 ( .A1(n16116), .A2(gray_img[505]), .B1(n15914), .B2(
        gray_img[1785]), .O(n17473) );
  AOI22S U23417 ( .A1(n17703), .A2(gray_img[633]), .B1(n17767), .B2(
        gray_img[1649]), .O(n17472) );
  AOI22S U23418 ( .A1(n17770), .A2(gray_img[497]), .B1(n15873), .B2(
        gray_img[2041]), .O(n17471) );
  INV1S U23419 ( .I(gray_img[881]), .O(n26375) );
  MOAI1S U23420 ( .A1(n17766), .A2(n26375), .B1(n17765), .B2(gray_img[1897]), 
        .O(n17470) );
  AN4B1S U23421 ( .I1(n17473), .I2(n17472), .I3(n17471), .B1(n17470), .O(
        n17491) );
  AOI22S U23422 ( .A1(n15913), .A2(gray_img[1505]), .B1(n17750), .B2(
        gray_img[481]), .O(n17477) );
  AOI22S U23423 ( .A1(n16000), .A2(gray_img[1121]), .B1(n17751), .B2(
        gray_img[1633]), .O(n17476) );
  AOI22S U23424 ( .A1(n15909), .A2(gray_img[225]), .B1(n15903), .B2(
        gray_img[1377]), .O(n17475) );
  MOAI1S U23425 ( .A1(n17753), .A2(intadd_4_CI), .B1(n17752), .B2(
        gray_img[353]), .O(n17474) );
  AN4B1S U23426 ( .I1(n17477), .I2(n17476), .I3(n17475), .B1(n17474), .O(
        n17490) );
  AOI22S U23427 ( .A1(n15902), .A2(gray_img[1761]), .B1(n17478), .B2(
        gray_img[97]), .O(n17482) );
  AOI22S U23428 ( .A1(n17758), .A2(gray_img[865]), .B1(n16165), .B2(
        gray_img[609]), .O(n17481) );
  AOI22S U23429 ( .A1(n17759), .A2(gray_img[1249]), .B1(n15901), .B2(
        gray_img[1889]), .O(n17480) );
  INV1S U23430 ( .I(gray_img[737]), .O(n26162) );
  MOAI1S U23431 ( .A1(n17760), .A2(n26162), .B1(n15900), .B2(gray_img[993]), 
        .O(n17479) );
  AN4B1S U23432 ( .I1(n17482), .I2(n17481), .I3(n17480), .B1(n17479), .O(
        n17489) );
  INV1S U23433 ( .I(gray_img[889]), .O(n26388) );
  MOAI1S U23434 ( .A1(n15946), .A2(n26388), .B1(n15911), .B2(gray_img[1913]), 
        .O(n17484) );
  MOAI1S U23435 ( .A1(n17745), .A2(intadd_103_CI), .B1(n15948), .B2(
        gray_img[1905]), .O(n17483) );
  NR2 U23436 ( .I1(n17484), .I2(n17483), .O(n17487) );
  AOI22S U23437 ( .A1(n15908), .A2(gray_img[1657]), .B1(n17743), .B2(
        gray_img[1641]), .O(n17486) );
  AOI22S U23438 ( .A1(n16137), .A2(gray_img[873]), .B1(n17744), .B2(
        gray_img[625]), .O(n17485) );
  ND3S U23439 ( .I1(n17487), .I2(n17486), .I3(n17485), .O(n17488) );
  AN4B1S U23440 ( .I1(n17491), .I2(n17490), .I3(n17489), .B1(n17488), .O(
        n17503) );
  AOI22S U23441 ( .A1(n15874), .A2(gray_img[1129]), .B1(n17804), .B2(
        gray_img[1401]), .O(n17495) );
  AOI22S U23442 ( .A1(n16001), .A2(gray_img[753]), .B1(n15875), .B2(
        gray_img[121]), .O(n17494) );
  AOI22S U23443 ( .A1(n17807), .A2(gray_img[1009]), .B1(n15951), .B2(
        gray_img[1265]), .O(n17493) );
  MOAI1S U23444 ( .A1(n17533), .A2(intadd_123_CI), .B1(n17805), .B2(
        gray_img[1769]), .O(n17492) );
  AN4B1S U23445 ( .I1(n17495), .I2(n17494), .I3(n17493), .B1(n17492), .O(
        n17501) );
  AOI22S U23446 ( .A1(n17796), .A2(gray_img[1385]), .B1(n17795), .B2(
        gray_img[1001]), .O(n17500) );
  AOI22S U23447 ( .A1(n15897), .A2(gray_img[2033]), .B1(n17797), .B2(
        gray_img[1513]), .O(n17499) );
  AOI22S U23448 ( .A1(n17605), .A2(gray_img[1137]), .B1(n15879), .B2(
        gray_img[1017]), .O(n17497) );
  AOI22S U23449 ( .A1(n17798), .A2(gray_img[369]), .B1(n15950), .B2(
        gray_img[241]), .O(n17496) );
  ND2S U23450 ( .I1(n17497), .I2(n17496), .O(n17498) );
  AN4B1S U23451 ( .I1(n17501), .I2(n17500), .I3(n17499), .B1(n17498), .O(
        n17502) );
  ND3S U23452 ( .I1(n17504), .I2(n17503), .I3(n17502), .O(n17554) );
  AOI22S U23453 ( .A1(n15908), .A2(gray_img[1561]), .B1(n17743), .B2(
        gray_img[1545]), .O(n17509) );
  AOI22S U23454 ( .A1(n15898), .A2(gray_img[793]), .B1(n15911), .B2(
        gray_img[1817]), .O(n17508) );
  AOI22S U23455 ( .A1(n15948), .A2(gray_img[1809]), .B1(n17709), .B2(
        gray_img[521]), .O(n17507) );
  INV1S U23456 ( .I(gray_img[529]), .O(n29051) );
  MOAI1S U23457 ( .A1(n17505), .A2(n29051), .B1(n16137), .B2(gray_img[777]), 
        .O(n17506) );
  AN4B1S U23458 ( .I1(n17509), .I2(n17508), .I3(n17507), .B1(n17506), .O(
        n17528) );
  AOI22S U23459 ( .A1(n16116), .A2(gray_img[409]), .B1(n15914), .B2(
        gray_img[1689]), .O(n17513) );
  AOI22S U23460 ( .A1(n17770), .A2(gray_img[401]), .B1(n15873), .B2(
        gray_img[1945]), .O(n17512) );
  AOI22S U23461 ( .A1(n15917), .A2(gray_img[785]), .B1(n17765), .B2(
        gray_img[1801]), .O(n17511) );
  INV1S U23462 ( .I(gray_img[537]), .O(n29063) );
  MOAI1S U23463 ( .A1(n17674), .A2(n29063), .B1(n17767), .B2(gray_img[1553]), 
        .O(n17510) );
  AN4B1S U23464 ( .I1(n17513), .I2(n17512), .I3(n17511), .B1(n17510), .O(
        n17527) );
  AOI22S U23465 ( .A1(n17752), .A2(gray_img[257]), .B1(n17696), .B2(
        gray_img[1921]), .O(n17517) );
  AOI22S U23466 ( .A1(n15913), .A2(gray_img[1409]), .B1(n17750), .B2(
        gray_img[385]), .O(n17516) );
  AOI22S U23467 ( .A1(n15909), .A2(gray_img[129]), .B1(n15903), .B2(
        gray_img[1281]), .O(n17515) );
  INV1S U23468 ( .I(gray_img[1537]), .O(n26588) );
  MOAI1S U23469 ( .A1(n15942), .A2(n26588), .B1(n16000), .B2(gray_img[1025]), 
        .O(n17514) );
  AN4B1S U23470 ( .I1(n17517), .I2(n17516), .I3(n17515), .B1(n17514), .O(
        n17526) );
  MOAI1S U23471 ( .A1(n17640), .A2(intadd_8_CI), .B1(n17758), .B2(
        gray_img[769]), .O(n17520) );
  MOAI1S U23472 ( .A1(n17518), .A2(intadd_88_CI), .B1(n15901), .B2(
        gray_img[1793]), .O(n17519) );
  NR2 U23473 ( .I1(n17520), .I2(n17519), .O(n17524) );
  AOI22S U23474 ( .A1(n15900), .A2(gray_img[897]), .B1(n17639), .B2(
        gray_img[641]), .O(n17523) );
  AOI22S U23475 ( .A1(n15902), .A2(gray_img[1665]), .B1(n15912), .B2(
        gray_img[1]), .O(n17522) );
  ND3S U23476 ( .I1(n17524), .I2(n17523), .I3(n17522), .O(n17525) );
  AN4B1S U23477 ( .I1(n17528), .I2(n17527), .I3(n17526), .B1(n17525), .O(
        n17552) );
  AOI22S U23478 ( .A1(n17778), .A2(gray_img[393]), .B1(n15895), .B2(
        gray_img[1433]), .O(n17532) );
  AOI22S U23479 ( .A1(n15877), .A2(gray_img[265]), .B1(n15899), .B2(
        gray_img[649]), .O(n17531) );
  AOI22S U23480 ( .A1(n15876), .A2(gray_img[1681]), .B1(n16188), .B2(
        gray_img[1177]), .O(n17530) );
  INV1S U23481 ( .I(gray_img[9]), .O(n23418) );
  MOAI1S U23482 ( .A1(n16002), .A2(n23418), .B1(n17591), .B2(gray_img[281]), 
        .O(n17529) );
  AN4B1S U23483 ( .I1(n17532), .I2(n17531), .I3(n17530), .B1(n17529), .O(
        n17550) );
  AOI22S U23484 ( .A1(n15874), .A2(gray_img[1033]), .B1(n17804), .B2(
        gray_img[1305]), .O(n17537) );
  AOI22S U23485 ( .A1(n16001), .A2(gray_img[657]), .B1(n15875), .B2(
        gray_img[25]), .O(n17536) );
  AOI22S U23486 ( .A1(n17807), .A2(gray_img[913]), .B1(n15951), .B2(
        gray_img[1169]), .O(n17535) );
  MOAI1S U23487 ( .A1(n17533), .A2(n27864), .B1(n17805), .B2(gray_img[1673]), 
        .O(n17534) );
  AN4B1S U23488 ( .I1(n17537), .I2(n17536), .I3(n17535), .B1(n17534), .O(
        n17549) );
  AOI22S U23489 ( .A1(n15897), .A2(gray_img[1937]), .B1(n17797), .B2(
        gray_img[1417]), .O(n17541) );
  AOI22S U23490 ( .A1(n17605), .A2(gray_img[1041]), .B1(n15879), .B2(
        gray_img[921]), .O(n17540) );
  AOI22S U23491 ( .A1(n17798), .A2(gray_img[273]), .B1(n15950), .B2(
        gray_img[145]), .O(n17539) );
  MOAI1S U23492 ( .A1(n17718), .A2(intadd_147_CI), .B1(n17796), .B2(
        gray_img[1289]), .O(n17538) );
  AN4B1S U23493 ( .I1(n17541), .I2(n17540), .I3(n17539), .B1(n17538), .O(
        n17548) );
  MOAI1S U23494 ( .A1(n15941), .A2(intadd_11_CI), .B1(n15949), .B2(
        gray_img[1425]), .O(n17543) );
  INV1S U23495 ( .I(gray_img[1297]), .O(n29747) );
  MOAI1S U23496 ( .A1(n15944), .A2(n29747), .B1(n17787), .B2(gray_img[137]), 
        .O(n17542) );
  NR2 U23497 ( .I1(n17543), .I2(n17542), .O(n17546) );
  AOI22S U23498 ( .A1(n15872), .A2(gray_img[1049]), .B1(n17785), .B2(
        gray_img[1161]), .O(n17545) );
  AOI22S U23499 ( .A1(n17786), .A2(gray_img[665]), .B1(n15866), .B2(
        gray_img[1929]), .O(n17544) );
  ND3S U23500 ( .I1(n17546), .I2(n17545), .I3(n17544), .O(n17547) );
  AN4B1S U23501 ( .I1(n17550), .I2(n17549), .I3(n17548), .B1(n17547), .O(
        n17551) );
  ND2S U23502 ( .I1(n17552), .I2(n17551), .O(n17553) );
  AOI22S U23503 ( .A1(n17554), .A2(n17819), .B1(n17553), .B2(n17688), .O(
        n17555) );
  NR2 U23504 ( .I1(n15996), .I2(n15870), .O(n17824) );
  FA1 U23505 ( .A(n17559), .B(n17558), .CI(n17557), .CO(n17572), .S(n17928) );
  FA1 U23506 ( .A(n17562), .B(n17561), .CI(n17560), .CO(n17571), .S(n17927) );
  NR2 U23507 ( .I1(n15996), .I2(n17868), .O(n17566) );
  NR2 U23508 ( .I1(n15992), .I2(n15871), .O(n17565) );
  HA1 U23509 ( .A(cro_mac[8]), .B(n17563), .C(n17557), .S(n17564) );
  NR2 U23510 ( .I1(n15994), .I2(n15943), .O(n17569) );
  NR2 U23511 ( .I1(n15997), .I2(n15870), .O(n17568) );
  NR2 U23512 ( .I1(n15992), .I2(n17957), .O(n17832) );
  NR2 U23513 ( .I1(n15994), .I2(n17873), .O(n17831) );
  NR2 U23514 ( .I1(n15993), .I2(n15943), .O(n17830) );
  NR2 U23515 ( .I1(n15991), .I2(n15871), .O(n17835) );
  NR2 U23516 ( .I1(n15995), .I2(n17868), .O(n17834) );
  NR2 U23517 ( .I1(n15995), .I2(n15870), .O(n17823) );
  FA1 U23518 ( .A(n17566), .B(n17565), .CI(n17564), .CO(n17932), .S(n17840) );
  FA1 U23519 ( .A(n17569), .B(n17568), .CI(n17567), .CO(n17931), .S(n17839) );
  NR2 U23520 ( .I1(n17940), .I2(n17942), .O(n17575) );
  FA1 U23521 ( .A(n17572), .B(n17571), .CI(n17570), .CO(n17963), .S(n17939) );
  INV1S U23522 ( .I(n17939), .O(n17574) );
  INV1S U23523 ( .I(n18007), .O(n17578) );
  ND2S U23524 ( .I1(n17577), .I2(n17576), .O(n18006) );
  ND2S U23525 ( .I1(n17578), .I2(n18006), .O(n17948) );
  NR2 U23526 ( .I1(n15991), .I2(n17957), .O(n17828) );
  NR2 U23527 ( .I1(n15994), .I2(n17868), .O(n17827) );
  NR2 U23528 ( .I1(n15994), .I2(n15870), .O(n17829) );
  AO222S U23529 ( .A1(template_reg[8]), .A2(n17581), .B1(template_reg[0]), 
        .B2(n17579), .C1(n17580), .C2(template_reg[16]), .O(n17590) );
  ND2S U23530 ( .I1(n17582), .I2(cnt_cro_3b3[0]), .O(n17588) );
  AOI22S U23531 ( .A1(n17584), .A2(template_reg[64]), .B1(n17583), .B2(
        template_reg[56]), .O(n17587) );
  ND2S U23532 ( .I1(n17585), .I2(template_reg[48]), .O(n17586) );
  NR2 U23533 ( .I1(n15990), .I2(n15871), .O(n17858) );
  AOI22S U23534 ( .A1(n17778), .A2(gray_img[456]), .B1(n15895), .B2(
        gray_img[1496]), .O(n17595) );
  AOI22S U23535 ( .A1(n15877), .A2(gray_img[328]), .B1(gray_img[712]), .B2(
        n15899), .O(n17594) );
  AOI22S U23536 ( .A1(n15876), .A2(gray_img[1744]), .B1(n16188), .B2(
        gray_img[1240]), .O(n17593) );
  MOAI1S U23537 ( .A1(n16002), .A2(intadd_130_A_0_), .B1(n17591), .B2(
        gray_img[344]), .O(n17592) );
  AN4B1S U23538 ( .I1(n17595), .I2(n17594), .I3(n17593), .B1(n17592), .O(
        n17615) );
  AOI22S U23539 ( .A1(n15874), .A2(gray_img[1096]), .B1(n17804), .B2(
        gray_img[1368]), .O(n17599) );
  AOI22S U23540 ( .A1(n17806), .A2(gray_img[216]), .B1(n17805), .B2(
        gray_img[1736]), .O(n17598) );
  AOI22S U23541 ( .A1(n17807), .A2(gray_img[976]), .B1(n15951), .B2(
        gray_img[1232]), .O(n17597) );
  MOAI1S U23542 ( .A1(n15868), .A2(intadd_188_A_0_), .B1(n16001), .B2(
        gray_img[720]), .O(n17596) );
  AN4B1S U23543 ( .I1(n17599), .I2(n17598), .I3(n17597), .B1(n17596), .O(
        n17614) );
  AOI22S U23544 ( .A1(n15872), .A2(gray_img[1112]), .B1(n17785), .B2(
        gray_img[1224]), .O(n17604) );
  AOI22S U23545 ( .A1(gray_img[1360]), .A2(n15878), .B1(n17787), .B2(
        gray_img[200]), .O(n17603) );
  AOI22S U23546 ( .A1(n17788), .A2(gray_img[80]), .B1(n15949), .B2(
        gray_img[1488]), .O(n17602) );
  INV1S U23547 ( .I(gray_img[1992]), .O(n17600) );
  MOAI1S U23548 ( .A1(n17600), .A2(n15894), .B1(n17786), .B2(gray_img[728]), 
        .O(n17601) );
  AN4B1S U23549 ( .I1(n17604), .I2(n17603), .I3(n17602), .B1(n17601), .O(
        n17613) );
  AOI22S U23550 ( .A1(gray_img[1104]), .A2(n17605), .B1(n15879), .B2(
        gray_img[984]), .O(n17608) );
  AOI22S U23551 ( .A1(n17606), .A2(gray_img[336]), .B1(n15950), .B2(
        gray_img[208]), .O(n17607) );
  AN2S U23552 ( .I1(n17608), .I2(n17607), .O(n17611) );
  AOI22S U23553 ( .A1(gray_img[1352]), .A2(n17796), .B1(n17795), .B2(
        gray_img[968]), .O(n17610) );
  AOI22S U23554 ( .A1(gray_img[2000]), .A2(n15897), .B1(n17797), .B2(
        gray_img[1480]), .O(n17609) );
  ND3S U23555 ( .I1(n17611), .I2(n17610), .I3(n17609), .O(n17612) );
  AN4B1S U23556 ( .I1(n17615), .I2(n17614), .I3(n17613), .B1(n17612), .O(
        n17638) );
  AOI22S U23557 ( .A1(n16116), .A2(gray_img[472]), .B1(gray_img[1752]), .B2(
        n15914), .O(n17619) );
  AOI22S U23558 ( .A1(n17770), .A2(gray_img[464]), .B1(n15873), .B2(
        gray_img[2008]), .O(n17618) );
  AOI22S U23559 ( .A1(n15917), .A2(gray_img[848]), .B1(n17765), .B2(
        gray_img[1864]), .O(n17617) );
  MOAI1S U23560 ( .A1(n17704), .A2(intadd_39_B_0_), .B1(n17703), .B2(
        gray_img[600]), .O(n17616) );
  AN4B1S U23561 ( .I1(n17619), .I2(n17618), .I3(n17617), .B1(n17616), .O(
        n17625) );
  AOI22S U23562 ( .A1(n15898), .A2(gray_img[856]), .B1(n15911), .B2(
        gray_img[1880]), .O(n17624) );
  AOI22S U23563 ( .A1(n15948), .A2(gray_img[1872]), .B1(n17709), .B2(
        gray_img[584]), .O(n17623) );
  AOI22S U23564 ( .A1(gray_img[1624]), .A2(n15908), .B1(n17743), .B2(
        gray_img[1608]), .O(n17621) );
  AOI22S U23565 ( .A1(n16137), .A2(gray_img[840]), .B1(n17744), .B2(
        gray_img[592]), .O(n17620) );
  ND2S U23566 ( .I1(n17621), .I2(n17620), .O(n17622) );
  AN4B1S U23567 ( .I1(n17625), .I2(n17624), .I3(n17623), .B1(n17622), .O(
        n17637) );
  AOI22S U23568 ( .A1(n15913), .A2(gray_img[1472]), .B1(n17750), .B2(
        gray_img[448]), .O(n17629) );
  AOI22S U23569 ( .A1(n16000), .A2(gray_img[1088]), .B1(gray_img[1600]), .B2(
        n17751), .O(n17628) );
  AOI22S U23570 ( .A1(n15909), .A2(gray_img[192]), .B1(n15903), .B2(
        gray_img[1344]), .O(n17627) );
  MOAI1S U23571 ( .A1(n17753), .A2(intadd_25_A_0_), .B1(n17752), .B2(
        gray_img[320]), .O(n17626) );
  AN4B1S U23572 ( .I1(n17629), .I2(n17628), .I3(n17627), .B1(n17626), .O(
        n17635) );
  AOI22S U23573 ( .A1(n15900), .A2(gray_img[960]), .B1(n17639), .B2(
        gray_img[704]), .O(n17634) );
  AOI22S U23574 ( .A1(n15902), .A2(gray_img[1728]), .B1(gray_img[64]), .B2(
        n15912), .O(n17633) );
  AOI22S U23575 ( .A1(n17758), .A2(gray_img[832]), .B1(n16165), .B2(
        gray_img[576]), .O(n17631) );
  AOI22S U23576 ( .A1(n17759), .A2(gray_img[1216]), .B1(n15901), .B2(
        gray_img[1856]), .O(n17630) );
  ND2S U23577 ( .I1(n17631), .I2(n17630), .O(n17632) );
  AN4B1S U23578 ( .I1(n17635), .I2(n17634), .I3(n17633), .B1(n17632), .O(
        n17636) );
  ND3S U23579 ( .I1(n17638), .I2(n17637), .I3(n17636), .O(n17691) );
  AOI22S U23580 ( .A1(gray_img[896]), .A2(n15900), .B1(n17639), .B2(
        gray_img[640]), .O(n17644) );
  AOI22S U23581 ( .A1(n15902), .A2(gray_img[1664]), .B1(n17478), .B2(
        gray_img[0]), .O(n17643) );
  AOI22S U23582 ( .A1(n17759), .A2(gray_img[1152]), .B1(gray_img[1792]), .B2(
        n15901), .O(n17642) );
  MOAI1S U23583 ( .A1(n17640), .A2(intadd_8_B_0_), .B1(n17758), .B2(
        gray_img[768]), .O(n17641) );
  AN4B1S U23584 ( .I1(n17644), .I2(n17643), .I3(n17642), .B1(n17641), .O(
        n17650) );
  AOI22S U23585 ( .A1(n15913), .A2(gray_img[1408]), .B1(gray_img[384]), .B2(
        n17750), .O(n17649) );
  AOI22S U23586 ( .A1(n16000), .A2(gray_img[1024]), .B1(gray_img[1536]), .B2(
        n17751), .O(n17648) );
  AOI22S U23587 ( .A1(gray_img[256]), .A2(n17752), .B1(n17696), .B2(
        gray_img[1920]), .O(n17646) );
  AOI22S U23588 ( .A1(n15909), .A2(gray_img[128]), .B1(n15903), .B2(
        gray_img[1280]), .O(n17645) );
  ND2S U23589 ( .I1(n17646), .I2(n17645), .O(n17647) );
  AN4B1S U23590 ( .I1(n17650), .I2(n17649), .I3(n17648), .B1(n17647), .O(
        n17687) );
  AOI22S U23591 ( .A1(n17778), .A2(gray_img[392]), .B1(gray_img[1432]), .B2(
        n15895), .O(n17654) );
  AOI22S U23592 ( .A1(n15877), .A2(gray_img[264]), .B1(n15899), .B2(
        gray_img[648]), .O(n17653) );
  AOI22S U23593 ( .A1(gray_img[1680]), .A2(n15876), .B1(n16188), .B2(
        gray_img[1176]), .O(n17652) );
  INV1S U23594 ( .I(gray_img[8]), .O(n22117) );
  MOAI1S U23595 ( .A1(n16002), .A2(n22117), .B1(n17780), .B2(gray_img[280]), 
        .O(n17651) );
  AN4B1S U23596 ( .I1(n17654), .I2(n17653), .I3(n17652), .B1(n17651), .O(
        n17673) );
  AOI22S U23597 ( .A1(gray_img[1936]), .A2(n15897), .B1(n17797), .B2(
        gray_img[1416]), .O(n17659) );
  AOI22S U23598 ( .A1(n17798), .A2(gray_img[272]), .B1(n15950), .B2(
        gray_img[144]), .O(n17658) );
  AOI22S U23599 ( .A1(gray_img[1040]), .A2(n17605), .B1(n15879), .B2(
        gray_img[920]), .O(n17657) );
  INV1S U23600 ( .I(gray_img[1288]), .O(n17655) );
  MOAI1S U23601 ( .A1(n17655), .A2(n15998), .B1(n17795), .B2(gray_img[904]), 
        .O(n17656) );
  AN4B1S U23602 ( .I1(n17659), .I2(n17658), .I3(n17657), .B1(n17656), .O(
        n17672) );
  AOI22S U23603 ( .A1(n17806), .A2(gray_img[152]), .B1(n17805), .B2(
        gray_img[1672]), .O(n17664) );
  AOI22S U23604 ( .A1(n16001), .A2(gray_img[656]), .B1(n15896), .B2(
        gray_img[24]), .O(n17663) );
  AOI22S U23605 ( .A1(n17807), .A2(gray_img[912]), .B1(n15951), .B2(
        gray_img[1168]), .O(n17662) );
  INV1S U23606 ( .I(gray_img[1304]), .O(n22102) );
  MOAI1S U23607 ( .A1(n17660), .A2(n22102), .B1(n15874), .B2(gray_img[1032]), 
        .O(n17661) );
  AN4B1S U23608 ( .I1(n17664), .I2(n17663), .I3(n17662), .B1(n17661), .O(
        n17671) );
  MOAI1S U23609 ( .A1(n15941), .A2(intadd_11_B_0_), .B1(n15949), .B2(
        gray_img[1424]), .O(n17666) );
  MOAI1S U23610 ( .A1(n15944), .A2(intadd_62_B_0_), .B1(n17787), .B2(
        gray_img[136]), .O(n17665) );
  NR2 U23611 ( .I1(n17666), .I2(n17665), .O(n17669) );
  AOI22S U23612 ( .A1(n15872), .A2(gray_img[1048]), .B1(n17785), .B2(
        gray_img[1160]), .O(n17668) );
  AOI22S U23613 ( .A1(gray_img[664]), .A2(n17786), .B1(n15866), .B2(
        gray_img[1928]), .O(n17667) );
  ND3S U23614 ( .I1(n17669), .I2(n17668), .I3(n17667), .O(n17670) );
  AN4B1S U23615 ( .I1(n17673), .I2(n17672), .I3(n17671), .B1(n17670), .O(
        n17686) );
  AOI22S U23616 ( .A1(n16116), .A2(gray_img[408]), .B1(n15914), .B2(
        gray_img[1688]), .O(n17678) );
  AOI22S U23617 ( .A1(gray_img[400]), .A2(n17770), .B1(n15873), .B2(
        gray_img[1944]), .O(n17677) );
  AOI22S U23618 ( .A1(n15917), .A2(gray_img[784]), .B1(n17765), .B2(
        gray_img[1800]), .O(n17676) );
  INV1S U23619 ( .I(gray_img[536]), .O(n29064) );
  MOAI1S U23620 ( .A1(n29064), .A2(n17674), .B1(n17767), .B2(gray_img[1552]), 
        .O(n17675) );
  AN4B1S U23621 ( .I1(n17678), .I2(n17677), .I3(n17676), .B1(n17675), .O(
        n17684) );
  AOI22S U23622 ( .A1(n15898), .A2(gray_img[792]), .B1(n15911), .B2(
        gray_img[1816]), .O(n17683) );
  AOI22S U23623 ( .A1(n15948), .A2(gray_img[1808]), .B1(n17709), .B2(
        gray_img[520]), .O(n17682) );
  AOI22S U23624 ( .A1(n15908), .A2(gray_img[1560]), .B1(n17743), .B2(
        gray_img[1544]), .O(n17680) );
  AOI22S U23625 ( .A1(n16137), .A2(gray_img[776]), .B1(n17744), .B2(
        gray_img[528]), .O(n17679) );
  ND2S U23626 ( .I1(n17680), .I2(n17679), .O(n17681) );
  AN4B1S U23627 ( .I1(n17684), .I2(n17683), .I3(n17682), .B1(n17681), .O(
        n17685) );
  ND3S U23628 ( .I1(n17687), .I2(n17686), .I3(n17685), .O(n17689) );
  AOI22S U23629 ( .A1(n17691), .A2(n17690), .B1(n17689), .B2(n17688), .O(
        n17822) );
  AOI22S U23630 ( .A1(n15902), .A2(gray_img[1760]), .B1(gray_img[96]), .B2(
        n15912), .O(n17695) );
  AOI22S U23631 ( .A1(n17758), .A2(gray_img[864]), .B1(n16165), .B2(
        gray_img[608]), .O(n17694) );
  AOI22S U23632 ( .A1(n17759), .A2(gray_img[1248]), .B1(n15901), .B2(
        gray_img[1888]), .O(n17693) );
  INV1S U23633 ( .I(gray_img[736]), .O(n26161) );
  MOAI1S U23634 ( .A1(n17760), .A2(n26161), .B1(n15900), .B2(gray_img[992]), 
        .O(n17692) );
  AN4B1S U23635 ( .I1(n17695), .I2(n17694), .I3(n17693), .B1(n17692), .O(
        n17702) );
  AOI22S U23636 ( .A1(n15913), .A2(gray_img[1504]), .B1(gray_img[480]), .B2(
        n17750), .O(n17701) );
  AOI22S U23637 ( .A1(n16000), .A2(gray_img[1120]), .B1(gray_img[1632]), .B2(
        n17751), .O(n17700) );
  AOI22S U23638 ( .A1(gray_img[352]), .A2(n17752), .B1(n17696), .B2(
        gray_img[2016]), .O(n17698) );
  AOI22S U23639 ( .A1(n15909), .A2(gray_img[224]), .B1(gray_img[1376]), .B2(
        n15903), .O(n17697) );
  ND2S U23640 ( .I1(n17698), .I2(n17697), .O(n17699) );
  AN4B1S U23641 ( .I1(n17702), .I2(n17701), .I3(n17700), .B1(n17699), .O(
        n17742) );
  AOI22S U23642 ( .A1(n16116), .A2(gray_img[504]), .B1(n15914), .B2(
        gray_img[1784]), .O(n17708) );
  AOI22S U23643 ( .A1(gray_img[496]), .A2(n17770), .B1(n15873), .B2(
        gray_img[2040]), .O(n17707) );
  AOI22S U23644 ( .A1(n15917), .A2(gray_img[880]), .B1(n17765), .B2(
        gray_img[1896]), .O(n17706) );
  INV1S U23645 ( .I(gray_img[1648]), .O(n22182) );
  MOAI1S U23646 ( .A1(n22182), .A2(n17704), .B1(n17703), .B2(gray_img[632]), 
        .O(n17705) );
  AN4B1S U23647 ( .I1(n17708), .I2(n17707), .I3(n17706), .B1(n17705), .O(
        n17715) );
  AOI22S U23648 ( .A1(n15898), .A2(gray_img[888]), .B1(gray_img[1912]), .B2(
        n15911), .O(n17714) );
  AOI22S U23649 ( .A1(n15948), .A2(gray_img[1904]), .B1(n17709), .B2(
        gray_img[616]), .O(n17713) );
  AOI22S U23650 ( .A1(n15908), .A2(gray_img[1656]), .B1(n17743), .B2(
        gray_img[1640]), .O(n17711) );
  AOI22S U23651 ( .A1(n16137), .A2(gray_img[872]), .B1(n17744), .B2(
        gray_img[624]), .O(n17710) );
  ND2S U23652 ( .I1(n17711), .I2(n17710), .O(n17712) );
  AN4B1S U23653 ( .I1(n17715), .I2(n17714), .I3(n17713), .B1(n17712), .O(
        n17741) );
  AOI22S U23654 ( .A1(n17716), .A2(gray_img[2032]), .B1(n17797), .B2(
        gray_img[1512]), .O(n17722) );
  AOI22S U23655 ( .A1(n17605), .A2(gray_img[1136]), .B1(n15879), .B2(
        gray_img[1016]), .O(n17721) );
  AOI22S U23656 ( .A1(n17717), .A2(gray_img[368]), .B1(n15950), .B2(
        gray_img[240]), .O(n17720) );
  INV1S U23657 ( .I(gray_img[1000]), .O(n22190) );
  MOAI1S U23658 ( .A1(n17718), .A2(n22190), .B1(n17796), .B2(gray_img[1384]), 
        .O(n17719) );
  AN4B1S U23659 ( .I1(n17722), .I2(n17721), .I3(n17720), .B1(n17719), .O(
        n17739) );
  AOI22S U23660 ( .A1(n16001), .A2(gray_img[752]), .B1(n15896), .B2(
        gray_img[120]), .O(n17727) );
  AOI22S U23661 ( .A1(n17807), .A2(gray_img[1008]), .B1(n15951), .B2(
        gray_img[1264]), .O(n17726) );
  AOI22S U23662 ( .A1(n15874), .A2(gray_img[1128]), .B1(n17804), .B2(
        gray_img[1400]), .O(n17725) );
  AOI22S U23663 ( .A1(n17806), .A2(gray_img[248]), .B1(n17805), .B2(
        gray_img[1768]), .O(n17724) );
  AN4S U23664 ( .I1(n17727), .I2(n17726), .I3(n17725), .I4(n17724), .O(n17738)
         );
  AOI22S U23665 ( .A1(n17778), .A2(gray_img[488]), .B1(n15895), .B2(
        gray_img[1528]), .O(n17731) );
  AOI22S U23666 ( .A1(gray_img[1776]), .A2(n15876), .B1(n16188), .B2(
        gray_img[1272]), .O(n17730) );
  AOI22S U23667 ( .A1(n17780), .A2(gray_img[376]), .B1(n17779), .B2(
        gray_img[104]), .O(n17729) );
  AOI22S U23668 ( .A1(n15877), .A2(gray_img[360]), .B1(gray_img[744]), .B2(
        n15899), .O(n17728) );
  AN4S U23669 ( .I1(n17731), .I2(n17730), .I3(n17729), .I4(n17728), .O(n17737)
         );
  AOI22S U23670 ( .A1(n15872), .A2(gray_img[1144]), .B1(n17785), .B2(
        gray_img[1256]), .O(n17735) );
  AOI22S U23671 ( .A1(gray_img[1392]), .A2(n15878), .B1(n17787), .B2(
        gray_img[232]), .O(n17734) );
  AOI22S U23672 ( .A1(n17788), .A2(gray_img[112]), .B1(n15949), .B2(
        gray_img[1520]), .O(n17733) );
  MOAI1S U23673 ( .A1(intadd_5_B_0_), .A2(n15894), .B1(n17786), .B2(
        gray_img[760]), .O(n17732) );
  AN4B1S U23674 ( .I1(n17735), .I2(n17734), .I3(n17733), .B1(n17732), .O(
        n17736) );
  AOI22S U23675 ( .A1(gray_img[1592]), .A2(n15908), .B1(n17743), .B2(
        gray_img[1576]), .O(n17749) );
  AOI22S U23676 ( .A1(n15898), .A2(gray_img[824]), .B1(n15911), .B2(
        gray_img[1848]), .O(n17748) );
  AOI22S U23677 ( .A1(n16137), .A2(gray_img[808]), .B1(n17744), .B2(
        gray_img[560]), .O(n17747) );
  MOAI1S U23678 ( .A1(n17745), .A2(intadd_137_A_0_), .B1(gray_img[1840]), .B2(
        n15948), .O(n17746) );
  AN4B1S U23679 ( .I1(n17749), .I2(n17748), .I3(n17747), .B1(n17746), .O(
        n17777) );
  AOI22S U23680 ( .A1(n15913), .A2(gray_img[1440]), .B1(n17750), .B2(
        gray_img[416]), .O(n17757) );
  AOI22S U23681 ( .A1(n16000), .A2(gray_img[1056]), .B1(gray_img[1568]), .B2(
        n17751), .O(n17756) );
  AOI22S U23682 ( .A1(n15909), .A2(gray_img[160]), .B1(gray_img[1312]), .B2(
        n15903), .O(n17755) );
  MOAI1S U23683 ( .A1(n17753), .A2(intadd_28_A_0_), .B1(n17752), .B2(
        gray_img[288]), .O(n17754) );
  AN4B1S U23684 ( .I1(n17757), .I2(n17756), .I3(n17755), .B1(n17754), .O(
        n17776) );
  AOI22S U23685 ( .A1(n15902), .A2(gray_img[1696]), .B1(n15912), .B2(
        gray_img[32]), .O(n17764) );
  AOI22S U23686 ( .A1(n17758), .A2(gray_img[800]), .B1(gray_img[544]), .B2(
        n16165), .O(n17763) );
  AOI22S U23687 ( .A1(n17759), .A2(gray_img[1184]), .B1(n15901), .B2(
        gray_img[1824]), .O(n17762) );
  INV1S U23688 ( .I(gray_img[672]), .O(n22046) );
  MOAI1S U23689 ( .A1(n17760), .A2(n22046), .B1(n15900), .B2(gray_img[928]), 
        .O(n17761) );
  AN4B1S U23690 ( .I1(n17764), .I2(n17763), .I3(n17762), .B1(n17761), .O(
        n17775) );
  INV1S U23691 ( .I(gray_img[816]), .O(n26097) );
  MOAI1S U23692 ( .A1(n17766), .A2(n26097), .B1(n17765), .B2(gray_img[1832]), 
        .O(n17769) );
  MOAI1S U23693 ( .A1(n17674), .A2(intadd_189_B_0_), .B1(n17767), .B2(
        gray_img[1584]), .O(n17768) );
  NR2 U23694 ( .I1(n17769), .I2(n17768), .O(n17773) );
  AOI22S U23695 ( .A1(n16116), .A2(gray_img[440]), .B1(gray_img[1720]), .B2(
        n15914), .O(n17772) );
  AOI22S U23696 ( .A1(gray_img[432]), .A2(n17770), .B1(n15873), .B2(
        gray_img[1976]), .O(n17771) );
  ND3S U23697 ( .I1(n17773), .I2(n17772), .I3(n17771), .O(n17774) );
  AN4B1S U23698 ( .I1(n17777), .I2(n17776), .I3(n17775), .B1(n17774), .O(
        n17816) );
  AOI22S U23699 ( .A1(n17778), .A2(gray_img[424]), .B1(gray_img[1464]), .B2(
        n15895), .O(n17784) );
  AOI22S U23700 ( .A1(n17780), .A2(gray_img[312]), .B1(gray_img[40]), .B2(
        n17779), .O(n17783) );
  AOI22S U23701 ( .A1(n15876), .A2(gray_img[1712]), .B1(n16188), .B2(
        gray_img[1208]), .O(n17782) );
  MOAI1S U23702 ( .A1(n16518), .A2(intadd_16_B_0_), .B1(n15899), .B2(
        gray_img[680]), .O(n17781) );
  AN4B1S U23703 ( .I1(n17784), .I2(n17783), .I3(n17782), .B1(n17781), .O(
        n17794) );
  AOI22S U23704 ( .A1(n15872), .A2(gray_img[1080]), .B1(gray_img[1192]), .B2(
        n17785), .O(n17793) );
  AOI22S U23705 ( .A1(n17786), .A2(gray_img[696]), .B1(n15866), .B2(
        gray_img[1960]), .O(n17792) );
  AOI22S U23706 ( .A1(n15878), .A2(gray_img[1328]), .B1(n17787), .B2(
        gray_img[168]), .O(n17790) );
  AOI22S U23707 ( .A1(n17788), .A2(gray_img[48]), .B1(n15949), .B2(
        gray_img[1456]), .O(n17789) );
  ND2S U23708 ( .I1(n17790), .I2(n17789), .O(n17791) );
  AN4B1S U23709 ( .I1(n17794), .I2(n17793), .I3(n17792), .B1(n17791), .O(
        n17815) );
  AOI22S U23710 ( .A1(n17796), .A2(gray_img[1320]), .B1(n17795), .B2(
        gray_img[936]), .O(n17803) );
  AOI22S U23711 ( .A1(gray_img[1968]), .A2(n15897), .B1(n17797), .B2(
        gray_img[1448]), .O(n17802) );
  AOI22S U23712 ( .A1(gray_img[1072]), .A2(n17605), .B1(n15879), .B2(
        gray_img[952]), .O(n17801) );
  INV1S U23713 ( .I(n17798), .O(n17799) );
  MOAI1S U23714 ( .A1(n17799), .A2(intadd_14_CI), .B1(n15950), .B2(
        gray_img[176]), .O(n17800) );
  AN4B1S U23715 ( .I1(n17803), .I2(n17802), .I3(n17801), .B1(n17800), .O(
        n17813) );
  AOI22S U23716 ( .A1(gray_img[688]), .A2(n16001), .B1(n15896), .B2(
        gray_img[56]), .O(n17812) );
  AOI22S U23717 ( .A1(n17723), .A2(gray_img[1064]), .B1(gray_img[1336]), .B2(
        n17804), .O(n17811) );
  AOI22S U23718 ( .A1(n17806), .A2(gray_img[184]), .B1(n17805), .B2(
        gray_img[1704]), .O(n17809) );
  AOI22S U23719 ( .A1(n17807), .A2(gray_img[944]), .B1(n15951), .B2(
        gray_img[1200]), .O(n17808) );
  ND2S U23720 ( .I1(n17809), .I2(n17808), .O(n17810) );
  AN4B1S U23721 ( .I1(n17813), .I2(n17812), .I3(n17811), .B1(n17810), .O(
        n17814) );
  ND3S U23722 ( .I1(n17816), .I2(n17815), .I3(n17814), .O(n17818) );
  AOI22S U23723 ( .A1(n17820), .A2(n17819), .B1(n17818), .B2(n17817), .O(
        n17821) );
  NR2 U23724 ( .I1(n15996), .I2(n15945), .O(n17857) );
  HA1 U23725 ( .A(cro_mac[6]), .B(n17823), .C(n17833), .S(n17856) );
  XNR2HS U23726 ( .I1(n17852), .I2(n17851), .O(n17825) );
  NR2 U23727 ( .I1(n15990), .I2(n17973), .O(n17850) );
  NR2 U23728 ( .I1(n15997), .I2(n15945), .O(n17849) );
  HA1 U23729 ( .A(cro_mac[7]), .B(n17824), .C(n17845), .S(n17848) );
  XNR2HS U23730 ( .I1(n17825), .I2(n17853), .O(n17867) );
  FA1 U23731 ( .A(n17828), .B(n17827), .CI(n17826), .CO(n17852), .S(n17864) );
  NR2 U23732 ( .I1(n15990), .I2(n17957), .O(n17900) );
  NR2 U23733 ( .I1(n15995), .I2(n15945), .O(n17899) );
  HA1 U23734 ( .A(cro_mac[5]), .B(n17829), .C(n17826), .S(n17898) );
  NR2 U23735 ( .I1(n15992), .I2(n15943), .O(n17838) );
  NR2 U23736 ( .I1(n15993), .I2(n17873), .O(n17837) );
  NR2 U23737 ( .I1(n15991), .I2(n15943), .O(n17861) );
  NR2 U23738 ( .I1(n15993), .I2(n17868), .O(n17860) );
  NR2 U23739 ( .I1(n15993), .I2(n15870), .O(n17872) );
  FA1 U23740 ( .A(n17832), .B(n17831), .CI(n17830), .CO(n17567), .S(n17844) );
  FA1 U23741 ( .A(n17835), .B(n17834), .CI(n17833), .CO(n17841), .S(n17843) );
  FA1 U23742 ( .A(n17838), .B(n17837), .CI(n17836), .CO(n17842), .S(n17862) );
  FA1 U23743 ( .A(n17841), .B(n17840), .CI(n17839), .CO(n17930), .S(n17926) );
  FA1 U23744 ( .A(n17844), .B(n17843), .CI(n17842), .CO(n17925), .S(n17865) );
  FA1 U23745 ( .A(n17847), .B(n17846), .CI(n17845), .CO(n17929), .S(n17935) );
  FA1 U23746 ( .A(n17850), .B(n17849), .CI(n17848), .CO(n17934), .S(n17853) );
  NR2 U23747 ( .I1(n17852), .I2(n17853), .O(n17855) );
  NR2 U23748 ( .I1(n17920), .I2(n17921), .O(n30167) );
  FA1 U23749 ( .A(n17858), .B(n17857), .CI(n17856), .CO(n17851), .S(n17915) );
  NR2 U23750 ( .I1(n15992), .I2(n17873), .O(n17897) );
  NR2 U23751 ( .I1(n15991), .I2(n17873), .O(n17871) );
  NR2 U23752 ( .I1(n15992), .I2(n17868), .O(n17870) );
  NR2 U23753 ( .I1(n15992), .I2(n15870), .O(n17874) );
  FA1 U23754 ( .A(n17861), .B(n17860), .CI(n17859), .CO(n17836), .S(n17895) );
  FA1 U23755 ( .A(n17864), .B(n17863), .CI(n17862), .CO(n17866), .S(n17913) );
  FA1 U23756 ( .A(n17867), .B(n17866), .CI(n17865), .CO(n17920), .S(n17919) );
  NR2 U23757 ( .I1(n17918), .I2(n17919), .O(n30175) );
  NR2 U23758 ( .I1(n30167), .I2(n30175), .O(n17923) );
  NR2 U23759 ( .I1(n15991), .I2(n17868), .O(n17880) );
  NR2 U23760 ( .I1(n15990), .I2(n17868), .O(n17881) );
  NR2 U23761 ( .I1(n15991), .I2(n15870), .O(n17884) );
  NR2 U23762 ( .I1(n15992), .I2(n15945), .O(n17883) );
  NR2 U23763 ( .I1(n15990), .I2(n15870), .O(n17885) );
  FA1 U23764 ( .A(n17871), .B(n17870), .CI(n17869), .CO(n17896), .S(n17906) );
  NR2 U23765 ( .I1(n15990), .I2(n15943), .O(n17903) );
  NR2 U23766 ( .I1(n15994), .I2(n15945), .O(n17902) );
  HA1 U23767 ( .A(cro_mac[4]), .B(n17872), .C(n17859), .S(n17901) );
  NR2 U23768 ( .I1(n15990), .I2(n17873), .O(n17877) );
  NR2 U23769 ( .I1(n15993), .I2(n15945), .O(n17876) );
  HA1 U23770 ( .A(cro_mac[3]), .B(n17874), .C(n17869), .S(n17875) );
  NR2 U23771 ( .I1(n17893), .I2(n17894), .O(n30193) );
  FA1 U23772 ( .A(n17877), .B(n17876), .CI(n17875), .CO(n17904), .S(n17891) );
  FA1 U23773 ( .A(n17880), .B(n17879), .CI(n17878), .CO(n17893), .S(n17892) );
  NR2 U23774 ( .I1(n17891), .I2(n17892), .O(n30199) );
  FA1 U23775 ( .A(n17884), .B(n17883), .CI(n17882), .CO(n17878), .S(n17889) );
  NR2 U23776 ( .I1(n15991), .I2(n15945), .O(n17886) );
  NR2 U23777 ( .I1(n17886), .I2(n17887), .O(n30210) );
  NR2 U23778 ( .I1(n15990), .I2(n15945), .O(n30215) );
  ND2S U23779 ( .I1(n30215), .I2(cro_mac[0]), .O(n30216) );
  ND2S U23780 ( .I1(n17887), .I2(n17886), .O(n30211) );
  OAI12HS U23781 ( .B1(n30210), .B2(n30216), .A1(n30211), .O(n30208) );
  ND2S U23782 ( .I1(n17889), .I2(n17888), .O(n30205) );
  INV1S U23783 ( .I(n30205), .O(n17890) );
  AOI12HS U23784 ( .B1(n30206), .B2(n30208), .A1(n17890), .O(n30203) );
  ND2S U23785 ( .I1(n17892), .I2(n17891), .O(n30200) );
  ND2S U23786 ( .I1(n17894), .I2(n17893), .O(n30194) );
  OAI12HS U23787 ( .B1(n30193), .B2(n30197), .A1(n30194), .O(n30190) );
  FA1 U23788 ( .A(n17900), .B(n17899), .CI(n17898), .CO(n17863), .S(n17912) );
  FA1 U23789 ( .A(n17903), .B(n17902), .CI(n17901), .CO(n17911), .S(n17905) );
  OR2 U23790 ( .I1(n17907), .I2(n17908), .O(n30189) );
  ND2S U23791 ( .I1(n17908), .I2(n17907), .O(n30188) );
  INV1S U23792 ( .I(n30188), .O(n17909) );
  AOI12HS U23793 ( .B1(n30190), .B2(n30189), .A1(n17909), .O(n30186) );
  FA1 U23794 ( .A(n17915), .B(n17914), .CI(n17913), .CO(n17918), .S(n17917) );
  NR2 U23795 ( .I1(n17916), .I2(n17917), .O(n30182) );
  ND2S U23796 ( .I1(n17917), .I2(n17916), .O(n30183) );
  OAI12HS U23797 ( .B1(n30186), .B2(n30182), .A1(n30183), .O(n30170) );
  ND2S U23798 ( .I1(n17919), .I2(n17918), .O(n30176) );
  ND2S U23799 ( .I1(n17921), .I2(n17920), .O(n30168) );
  OAI12HS U23800 ( .B1(n30167), .B2(n30176), .A1(n30168), .O(n17922) );
  INV2 U23801 ( .I(n17972), .O(n30163) );
  FA1 U23802 ( .A(n17926), .B(n17925), .CI(n17924), .CO(n17943), .S(n17921) );
  FA1 U23803 ( .A(n17929), .B(n17928), .CI(n17927), .CO(n17940), .S(n17938) );
  FA1 U23804 ( .A(n17932), .B(n17931), .CI(n17930), .CO(n17942), .S(n17937) );
  FA1 U23805 ( .A(n17935), .B(n17934), .CI(n17933), .CO(n17936), .S(n17924) );
  NR2 U23806 ( .I1(n17943), .I2(n17944), .O(n30155) );
  FA1 U23807 ( .A(n17938), .B(n17937), .CI(n17936), .CO(n17945), .S(n17944) );
  XNR2HS U23808 ( .I1(n17940), .I2(n17939), .O(n17941) );
  NR2 U23809 ( .I1(n17945), .I2(n17946), .O(n30152) );
  NR2 U23810 ( .I1(n30155), .I2(n30152), .O(n18003) );
  ND2S U23811 ( .I1(n17944), .I2(n17943), .O(n30161) );
  ND2S U23812 ( .I1(n17946), .I2(n17945), .O(n30153) );
  OAI12HS U23813 ( .B1(n30152), .B2(n30161), .A1(n30153), .O(n18005) );
  AOI12HS U23814 ( .B1(n30163), .B2(n18003), .A1(n18005), .O(n17947) );
  XOR2HS U23815 ( .I1(n17948), .I2(n17947), .O(n17952) );
  INV1S U23816 ( .I(n17949), .O(n17951) );
  NR2 U23817 ( .I1(n17951), .I2(n17950), .O(n30218) );
  MOAI1 U23818 ( .A1(n30220), .A2(n17953), .B1(n17952), .B2(n30218), .O(n13600) );
  INV1S U23819 ( .I(cro_mac[17]), .O(n18017) );
  FA1 U23820 ( .A(n17956), .B(n17955), .CI(n17954), .CO(n17986), .S(n17960) );
  NR2 U23821 ( .I1(n15997), .I2(n17957), .O(n17980) );
  NR2 U23822 ( .I1(n15995), .I2(n17973), .O(n17975) );
  NR2 U23823 ( .I1(n15996), .I2(n15871), .O(n17974) );
  FA1 U23824 ( .A(n17962), .B(n17961), .CI(n17960), .CO(n17984), .S(n17964) );
  FA1 U23825 ( .A(n17965), .B(n17964), .CI(n17963), .CO(n17967), .S(n17576) );
  NR2 U23826 ( .I1(n17966), .I2(n17967), .O(n18000) );
  NR2 U23827 ( .I1(n18000), .I2(n18007), .O(n17969) );
  ND2P U23828 ( .I1(n18003), .I2(n17969), .O(n17971) );
  ND2S U23829 ( .I1(n17967), .I2(n17966), .O(n18001) );
  OAI12HS U23830 ( .B1(n18000), .B2(n18006), .A1(n18001), .O(n17968) );
  AOI12H U23831 ( .B1(n18005), .B2(n17969), .A1(n17968), .O(n17970) );
  OAI12HP U23832 ( .B1(n17972), .B2(n17971), .A1(n17970), .O(n30148) );
  NR2 U23833 ( .I1(n15997), .I2(n17973), .O(n17988) );
  NR2 U23834 ( .I1(n15996), .I2(n17973), .O(n17977) );
  NR2 U23835 ( .I1(n15997), .I2(n15871), .O(n17976) );
  FA1S U23836 ( .A(cro_mac[13]), .B(n17977), .CI(n17976), .CO(n17987), .S(
        n17982) );
  FA1 U23837 ( .A(n17980), .B(n17979), .CI(n17978), .CO(n17981), .S(n17985) );
  NR2 U23838 ( .I1(n17991), .I2(n17992), .O(n18046) );
  NR2 U23839 ( .I1(n17989), .I2(n17990), .O(n18049) );
  NR2 U23840 ( .I1(n18046), .I2(n18049), .O(n18041) );
  INV1S U23841 ( .I(cro_mac[16]), .O(n18035) );
  FA1S U23842 ( .A(cro_mac[14]), .B(n17988), .CI(n17987), .CO(n17993), .S(
        n17991) );
  NR2 U23843 ( .I1(cro_mac[15]), .I2(n17993), .O(n18037) );
  NR2 U23844 ( .I1(n18035), .I2(n18037), .O(n17995) );
  ND2S U23845 ( .I1(n18041), .I2(n17995), .O(n18015) );
  INV1S U23846 ( .I(n18015), .O(n17997) );
  ND2S U23847 ( .I1(n17990), .I2(n17989), .O(n30146) );
  OAI12HS U23848 ( .B1(n30146), .B2(n18046), .A1(n18047), .O(n18040) );
  NR2 U23849 ( .I1(n18035), .I2(n18038), .O(n17994) );
  AOI12HS U23850 ( .B1(n18040), .B2(n17995), .A1(n17994), .O(n18016) );
  INV1S U23851 ( .I(n18016), .O(n17996) );
  AOI12HS U23852 ( .B1(n30148), .B2(n17997), .A1(n17996), .O(n17998) );
  XOR2HS U23853 ( .I1(n18017), .I2(n17998), .O(n17999) );
  MOAI1 U23854 ( .A1(n30220), .A2(n18017), .B1(n17999), .B2(n30218), .O(n13594) );
  INV1S U23855 ( .I(cro_mac[12]), .O(n18014) );
  INV1S U23856 ( .I(n18000), .O(n18002) );
  INV1S U23857 ( .I(n18003), .O(n18004) );
  NR2 U23858 ( .I1(n18007), .I2(n18004), .O(n18010) );
  INV1S U23859 ( .I(n18005), .O(n18008) );
  OAI12HS U23860 ( .B1(n18008), .B2(n18007), .A1(n18006), .O(n18009) );
  AOI12HS U23861 ( .B1(n18010), .B2(n30163), .A1(n18009), .O(n18011) );
  XOR2HS U23862 ( .I1(n18012), .I2(n18011), .O(n18013) );
  MOAI1 U23863 ( .A1(n30220), .A2(n18014), .B1(n18013), .B2(n30218), .O(n13599) );
  INV1S U23864 ( .I(cro_mac[18]), .O(n18019) );
  NR2 U23865 ( .I1(n18017), .I2(n18015), .O(n18021) );
  NR2 U23866 ( .I1(n18017), .I2(n18016), .O(n18023) );
  AOI12HS U23867 ( .B1(n30148), .B2(n18021), .A1(n18023), .O(n18018) );
  XOR2HS U23868 ( .I1(n18019), .I2(n18018), .O(n18020) );
  MOAI1 U23869 ( .A1(n30220), .A2(n18019), .B1(n18020), .B2(n30218), .O(n13593) );
  INV1S U23870 ( .I(cro_mac[19]), .O(n18028) );
  ND2S U23871 ( .I1(n18021), .I2(cro_mac[18]), .O(n18022) );
  INV1S U23872 ( .I(n18022), .O(n18026) );
  ND2S U23873 ( .I1(n18023), .I2(cro_mac[18]), .O(n18024) );
  INV1S U23874 ( .I(n18024), .O(n18025) );
  AOI12HS U23875 ( .B1(n30148), .B2(n18026), .A1(n18025), .O(n18027) );
  XOR2HS U23876 ( .I1(n18028), .I2(n18027), .O(n18029) );
  MOAI1 U23877 ( .A1(n30220), .A2(n18028), .B1(n18029), .B2(n30218), .O(n13592) );
  INV1S U23878 ( .I(n18041), .O(n18030) );
  NR2 U23879 ( .I1(n18037), .I2(n18030), .O(n18033) );
  INV1S U23880 ( .I(n18040), .O(n18031) );
  OAI12HS U23881 ( .B1(n18031), .B2(n18037), .A1(n18038), .O(n18032) );
  AOI12HS U23882 ( .B1(n30148), .B2(n18033), .A1(n18032), .O(n18034) );
  XOR2HS U23883 ( .I1(n18035), .I2(n18034), .O(n18036) );
  MOAI1 U23884 ( .A1(n30220), .A2(n18035), .B1(n18036), .B2(n30218), .O(n13595) );
  INV1S U23885 ( .I(cro_mac[15]), .O(n18045) );
  INV1S U23886 ( .I(n18037), .O(n18039) );
  ND2S U23887 ( .I1(n18039), .I2(n18038), .O(n18043) );
  AOI12HS U23888 ( .B1(n30148), .B2(n18041), .A1(n18040), .O(n18042) );
  XOR2HS U23889 ( .I1(n18043), .I2(n18042), .O(n18044) );
  MOAI1 U23890 ( .A1(n30220), .A2(n18045), .B1(n18044), .B2(n30218), .O(n13596) );
  INV1S U23891 ( .I(cro_mac[14]), .O(n18054) );
  INV1S U23892 ( .I(n18046), .O(n18048) );
  INV1S U23893 ( .I(n18049), .O(n30147) );
  INV1S U23894 ( .I(n30146), .O(n18050) );
  AOI12HS U23895 ( .B1(n30148), .B2(n30147), .A1(n18050), .O(n18051) );
  XOR2HS U23896 ( .I1(n18052), .I2(n18051), .O(n18053) );
  MOAI1 U23897 ( .A1(n30220), .A2(n18054), .B1(n18053), .B2(n30218), .O(n13597) );
  INV1S U23898 ( .I(image[7]), .O(n30423) );
  NR2P U23899 ( .I1(cnt_dyn[0]), .I2(n30349), .O(n30451) );
  INV2 U23900 ( .I(n30451), .O(n30452) );
  MOAI1S U23901 ( .A1(n30423), .A2(n30452), .B1(n18055), .B2(n30349), .O(
        n15823) );
  INV1S U23902 ( .I(gray_img[1471]), .O(n21934) );
  INV1S U23903 ( .I(gray_img[1469]), .O(n18062) );
  INV1S U23904 ( .I(gray_img[1468]), .O(n18060) );
  INV1S U23905 ( .I(gray_img[1467]), .O(n18058) );
  INV1S U23906 ( .I(gray_img[1466]), .O(n22380) );
  FA1S U23907 ( .A(gray_img[1337]), .B(gray_img[1336]), .CI(intadd_134_CI), 
        .CO(n18056) );
  FA1S U23908 ( .A(n22380), .B(gray_img[1338]), .CI(n18056), .CO(n18057) );
  FA1S U23909 ( .A(n18058), .B(gray_img[1339]), .CI(n18057), .CO(n18059) );
  FA1S U23910 ( .A(n18060), .B(gray_img[1340]), .CI(n18059), .CO(n18061) );
  MXL2HS U23911 ( .A(gray_img[1470]), .B(gray_img[1342]), .S(n29341), .OB(
        n18101) );
  INV1S U23912 ( .I(gray_img[1335]), .O(n18066) );
  INV1S U23913 ( .I(gray_img[1463]), .O(n18081) );
  ND2S U23914 ( .I1(n18066), .I2(n18081), .O(n25311) );
  NR2 U23915 ( .I1(gray_img[1471]), .I2(gray_img[1343]), .O(n25312) );
  INV1S U23916 ( .I(gray_img[1462]), .O(n18080) );
  INV1S U23917 ( .I(gray_img[1461]), .O(n18075) );
  INV1S U23918 ( .I(gray_img[1460]), .O(n18073) );
  INV1S U23919 ( .I(gray_img[1459]), .O(n18071) );
  INV1S U23920 ( .I(gray_img[1458]), .O(n18069) );
  INV1S U23921 ( .I(gray_img[1457]), .O(n18067) );
  FA1S U23922 ( .A(gray_img[1329]), .B(gray_img[1328]), .CI(n18067), .CO(
        n18068) );
  FA1S U23923 ( .A(n18069), .B(gray_img[1330]), .CI(n18068), .CO(n18070) );
  FA1S U23924 ( .A(n18071), .B(gray_img[1331]), .CI(n18070), .CO(n18072) );
  INV1S U23925 ( .I(gray_img[1333]), .O(n18077) );
  INV1S U23926 ( .I(gray_img[1334]), .O(n18076) );
  AOI22S U23927 ( .A1(n18077), .A2(gray_img[1461]), .B1(gray_img[1462]), .B2(
        n18076), .O(n18078) );
  AOI22S U23928 ( .A1(gray_img[1334]), .A2(n18080), .B1(n18079), .B2(n18078), 
        .O(n18083) );
  NR2 U23929 ( .I1(gray_img[1335]), .I2(n18081), .O(n18082) );
  MXL2HS U23930 ( .A(gray_img[1469]), .B(gray_img[1341]), .S(n29341), .OB(
        n28897) );
  MXL2HS U23931 ( .A(gray_img[1468]), .B(gray_img[1340]), .S(n29341), .OB(
        n23205) );
  MXL2HS U23932 ( .A(gray_img[1467]), .B(gray_img[1339]), .S(n29341), .OB(
        n28907) );
  MXL2HS U23933 ( .A(gray_img[1466]), .B(gray_img[1338]), .S(n29341), .OB(
        n28912) );
  MXL2HS U23934 ( .A(gray_img[1465]), .B(gray_img[1337]), .S(n29341), .OB(
        n28917) );
  OR2 U23935 ( .I1(n29680), .I2(n18091), .O(n29340) );
  INV1S U23936 ( .I(n18091), .O(n18092) );
  INV1S U23937 ( .I(medfilt_cnt_d1[2]), .O(n18136) );
  NR2 U23938 ( .I1(n18819), .I2(n24972), .O(n25086) );
  NR2 U23939 ( .I1(n18537), .I2(n18532), .O(n25308) );
  INV1S U23940 ( .I(cnt_dyn_d1[2]), .O(n18138) );
  NR2 U23941 ( .I1(n18538), .I2(n18533), .O(n25340) );
  AOI22S U23942 ( .A1(n25086), .A2(n25308), .B1(n25085), .B2(n25340), .O(
        n18096) );
  OA12S U23943 ( .B1(gray_img[670]), .B2(n29427), .A1(n29344), .O(n18098) );
  MOAI1S U23944 ( .A1(n29344), .A2(gray_img[670]), .B1(n29825), .B2(n18098), 
        .O(n18099) );
  INV1S U23945 ( .I(gray_img[269]), .O(n18110) );
  INV1S U23946 ( .I(gray_img[396]), .O(n18107) );
  INV1S U23947 ( .I(gray_img[395]), .O(n18105) );
  INV1S U23948 ( .I(gray_img[394]), .O(n18103) );
  FA1S U23949 ( .A(gray_img[265]), .B(gray_img[264]), .CI(intadd_204_CI), .CO(
        n18102) );
  FA1S U23950 ( .A(n18103), .B(gray_img[266]), .CI(n18102), .CO(n18104) );
  INV1S U23951 ( .I(n18108), .O(n18109) );
  MXL2HS U23952 ( .A(gray_img[270]), .B(gray_img[398]), .S(n18126), .OB(n18144) );
  INV1S U23953 ( .I(gray_img[263]), .O(n18113) );
  INV1S U23954 ( .I(gray_img[391]), .O(n18125) );
  ND2S U23955 ( .I1(n18113), .I2(n18125), .O(n25319) );
  NR2 U23956 ( .I1(gray_img[271]), .I2(gray_img[399]), .O(n25320) );
  INV1S U23957 ( .I(gray_img[390]), .O(n18123) );
  INV1S U23958 ( .I(gray_img[389]), .O(n18121) );
  INV1S U23959 ( .I(gray_img[388]), .O(n18119) );
  INV1S U23960 ( .I(gray_img[387]), .O(n18117) );
  INV1S U23961 ( .I(gray_img[386]), .O(n18115) );
  MAO222S U23962 ( .A1(gray_img[256]), .B1(gray_img[257]), .C1(intadd_153_CI), 
        .O(n18114) );
  MAO222S U23963 ( .A1(n18115), .B1(gray_img[258]), .C1(n18114), .O(n18116) );
  FA1S U23964 ( .A(n18117), .B(gray_img[259]), .CI(n18116), .CO(n18118) );
  FA1S U23965 ( .A(n18119), .B(gray_img[260]), .CI(n18118), .CO(n18120) );
  MXL2HS U23966 ( .A(gray_img[269]), .B(gray_img[397]), .S(n18126), .OB(n30041) );
  MXL2HS U23967 ( .A(gray_img[268]), .B(gray_img[396]), .S(n18126), .OB(n30047) );
  MXL2HS U23968 ( .A(gray_img[267]), .B(gray_img[395]), .S(n18126), .OB(n30053) );
  MXL2HS U23969 ( .A(gray_img[266]), .B(gray_img[394]), .S(n18126), .OB(n30060) );
  MXL2HS U23970 ( .A(gray_img[264]), .B(gray_img[392]), .S(n18126), .OB(n23366) );
  MXL2HS U23971 ( .A(gray_img[265]), .B(gray_img[393]), .S(n18126), .OB(n30124) );
  MAO222 U23972 ( .A1(n23366), .B1(n30124), .C1(n30127), .O(n18127) );
  OR2 U23973 ( .I1(n29680), .I2(n18133), .O(n30125) );
  INV1S U23974 ( .I(n18133), .O(n18134) );
  NR2 U23975 ( .I1(n18883), .I2(n24997), .O(n25218) );
  NR2 U23976 ( .I1(n18509), .I2(n18537), .O(n25246) );
  NR2 U23977 ( .I1(n18510), .I2(n18538), .O(n25257) );
  AOI22S U23978 ( .A1(n25218), .A2(n25246), .B1(n25216), .B2(n25257), .O(
        n18140) );
  OA12S U23979 ( .B1(gray_img[134]), .B2(n29427), .A1(n30121), .O(n18141) );
  MOAI1S U23980 ( .A1(n30121), .A2(gray_img[134]), .B1(n29825), .B2(n18141), 
        .O(n18142) );
  BUF1 U23981 ( .I(rst_n), .O(n30454) );
  NR2 U23982 ( .I1(cs[2]), .I2(cs[0]), .O(n30388) );
  INV1S U23983 ( .I(n30388), .O(n18397) );
  NR2 U23984 ( .I1(n18145), .I2(n18397), .O(n24967) );
  INV1S U23985 ( .I(n24967), .O(n30391) );
  ND2S U23986 ( .I1(n25315), .I2(action_done), .O(n18148) );
  ND2S U23987 ( .I1(image_size_reg_set[1]), .I2(n30391), .O(n24900) );
  NR2 U23988 ( .I1(image_size_reg_set[0]), .I2(n18148), .O(n24899) );
  INV1S U23989 ( .I(n24899), .O(n18146) );
  MOAI1S U23990 ( .A1(n24900), .A2(n18146), .B1(image_size_reg_master[0]), 
        .B2(n24967), .O(n18147) );
  AO13S U23991 ( .B1(image_size_reg_set[0]), .B2(n30391), .B3(n18148), .A1(
        n18147), .O(n15756) );
  INV1S U23992 ( .I(cnt_bdyn[1]), .O(n30369) );
  INV1S U23993 ( .I(cnt_bdyn[0]), .O(n30372) );
  NR2 U23994 ( .I1(n30369), .I2(n30372), .O(n30302) );
  INV1S U23995 ( .I(cnt_bdyn[3]), .O(n30330) );
  NR2 U23996 ( .I1(n30364), .I2(n30330), .O(n21125) );
  INV1S U23997 ( .I(n21125), .O(n30361) );
  XOR2HS U23998 ( .I1(cnt_dyn_base[1]), .I2(cnt_dyn[1]), .O(n18151) );
  XOR2HS U23999 ( .I1(cnt_dyn_base[3]), .I2(cnt_dyn[3]), .O(n18150) );
  INV1S U24000 ( .I(cnt_dyn[2]), .O(n30305) );
  XNR2HS U24001 ( .I1(cnt_dyn_base[2]), .I2(n30305), .O(n18149) );
  NR3 U24002 ( .I1(n18151), .I2(n18150), .I3(n18149), .O(n18453) );
  XNR2HS U24003 ( .I1(cnt_dyn_base[0]), .I2(cnt_dyn[0]), .O(n18152) );
  NR2 U24004 ( .I1(n30361), .I2(n30359), .O(n18154) );
  ND2S U24005 ( .I1(cnt_bdyn[4]), .I2(n18154), .O(n18153) );
  INV1S U24006 ( .I(n18153), .O(n30356) );
  NR2 U24007 ( .I1(last_in_valid), .I2(n30387), .O(n30255) );
  ND2S U24008 ( .I1(cnt_bdyn[6]), .I2(n30358), .O(n30352) );
  OA112S U24009 ( .C1(cnt_bdyn[6]), .C2(n30358), .A1(n24942), .B1(n30352), .O(
        n15802) );
  OA112S U24010 ( .C1(cnt_bdyn[4]), .C2(n18154), .A1(n24942), .B1(n18153), .O(
        n15800) );
  OR2S U24011 ( .I1(cnt_dyn_base[1]), .I2(n24898), .O(n18167) );
  INV1S U24012 ( .I(cnt_dyn_base[3]), .O(n24903) );
  NR2 U24013 ( .I1(cnt_dyn_base[2]), .I2(n24903), .O(n18166) );
  INV1S U24014 ( .I(n18166), .O(n18177) );
  ND2S U24015 ( .I1(cnt_dyn_base[3]), .I2(cnt_dyn_base[2]), .O(n18173) );
  INV1S U24016 ( .I(cnt_dyn_base[1]), .O(n18398) );
  NR2 U24017 ( .I1(n18398), .I2(n24898), .O(n18375) );
  INV1S U24018 ( .I(n18375), .O(n18156) );
  AOI22S U24019 ( .A1(n18155), .A2(mem_data_out_reg_shift_0[75]), .B1(n18157), 
        .B2(mem_data_out_reg_shift_0[123]), .O(n18164) );
  INV1S U24020 ( .I(cnt_dyn_base[2]), .O(n24902) );
  NR2 U24021 ( .I1(cnt_dyn_base[3]), .I2(n24902), .O(n18160) );
  AN2 U24022 ( .I1(n18375), .I2(n18160), .O(n18360) );
  AOI22S U24023 ( .A1(n18158), .A2(mem_data_out_reg_shift_0[107]), .B1(n18360), 
        .B2(mem_data_out_reg_shift_0[59]), .O(n18163) );
  OR2S U24024 ( .I1(cnt_dyn_base[2]), .I2(cnt_dyn_base[3]), .O(n18175) );
  OR2S U24025 ( .I1(cnt_dyn_base[0]), .I2(n18398), .O(n18178) );
  INV1S U24026 ( .I(n18160), .O(n18181) );
  AOI22S U24027 ( .A1(n18159), .A2(mem_data_out_reg_shift_0[19]), .B1(n18161), 
        .B2(mem_data_out_reg_shift_0[51]), .O(n18162) );
  ND3S U24028 ( .I1(n18164), .I2(n18163), .I3(n18162), .O(n18188) );
  INV1S U24029 ( .I(n18385), .O(n18180) );
  NR2 U24030 ( .I1(cnt_dyn_base[2]), .I2(n18180), .O(n18383) );
  AN2S U24031 ( .I1(n18383), .I2(cnt_dyn_base[3]), .O(n18359) );
  ND2S U24032 ( .I1(n18359), .I2(mem_data_out_reg_shift_0[67]), .O(n18172) );
  AN2 U24033 ( .I1(n18375), .I2(n18166), .O(n18357) );
  AOI22S U24034 ( .A1(n18165), .A2(mem_data_out_reg_shift_0[43]), .B1(n18357), 
        .B2(mem_data_out_reg_shift_0[91]), .O(n18171) );
  AOI22S U24035 ( .A1(n18168), .A2(mem_data_out_reg_shift_0[11]), .B1(n18169), 
        .B2(mem_data_out_reg_shift_0[99]), .O(n18170) );
  ND3S U24036 ( .I1(n18172), .I2(n18171), .I3(n18170), .O(n18187) );
  ND2S U24037 ( .I1(n18392), .I2(mem_data_out_reg_shift_0[3]), .O(n18185) );
  INV1S U24038 ( .I(n18175), .O(n18176) );
  AN2 U24039 ( .I1(n18375), .I2(n18176), .O(n18358) );
  AOI22S U24040 ( .A1(n18174), .A2(mem_data_out_reg_shift_0[115]), .B1(n18358), 
        .B2(mem_data_out_reg_shift_0[27]), .O(n18184) );
  AOI22S U24041 ( .A1(n18179), .A2(mem_data_out_reg_shift_0[83]), .B1(n18182), 
        .B2(mem_data_out_reg_shift_0[35]), .O(n18183) );
  ND3S U24042 ( .I1(n18185), .I2(n18184), .I3(n18183), .O(n18186) );
  OR3S U24043 ( .I1(n18188), .I2(n18187), .I3(n18186), .O(n15829) );
  AOI22S U24044 ( .A1(n18155), .A2(mem_data_out_reg_shift_0[74]), .B1(n18157), 
        .B2(mem_data_out_reg_shift_0[122]), .O(n18191) );
  AOI22S U24045 ( .A1(n18158), .A2(mem_data_out_reg_shift_0[106]), .B1(n18360), 
        .B2(mem_data_out_reg_shift_0[58]), .O(n18190) );
  AOI22S U24046 ( .A1(n18159), .A2(mem_data_out_reg_shift_0[18]), .B1(n18161), 
        .B2(mem_data_out_reg_shift_0[50]), .O(n18189) );
  ND2S U24047 ( .I1(n18359), .I2(mem_data_out_reg_shift_0[66]), .O(n18194) );
  AOI22S U24048 ( .A1(n18165), .A2(mem_data_out_reg_shift_0[42]), .B1(n18357), 
        .B2(mem_data_out_reg_shift_0[90]), .O(n18193) );
  AOI22S U24049 ( .A1(n18168), .A2(mem_data_out_reg_shift_0[10]), .B1(n18169), 
        .B2(mem_data_out_reg_shift_0[98]), .O(n18192) );
  ND3S U24050 ( .I1(n18194), .I2(n18193), .I3(n18192), .O(n18199) );
  ND2S U24051 ( .I1(n18392), .I2(mem_data_out_reg_shift_0[2]), .O(n18197) );
  AOI22S U24052 ( .A1(n18174), .A2(mem_data_out_reg_shift_0[114]), .B1(n18358), 
        .B2(mem_data_out_reg_shift_0[26]), .O(n18196) );
  AOI22S U24053 ( .A1(n18179), .A2(mem_data_out_reg_shift_0[82]), .B1(n18182), 
        .B2(mem_data_out_reg_shift_0[34]), .O(n18195) );
  ND3S U24054 ( .I1(n18197), .I2(n18196), .I3(n18195), .O(n18198) );
  OR3S U24055 ( .I1(n18200), .I2(n18199), .I3(n18198), .O(n15830) );
  AOI22S U24056 ( .A1(n18155), .A2(mem_data_out_reg_shift_1[72]), .B1(n18157), 
        .B2(mem_data_out_reg_shift_1[120]), .O(n18203) );
  AOI22S U24057 ( .A1(n18158), .A2(mem_data_out_reg_shift_1[104]), .B1(n18360), 
        .B2(mem_data_out_reg_shift_1[56]), .O(n18202) );
  AOI22S U24058 ( .A1(n18159), .A2(mem_data_out_reg_shift_1[16]), .B1(n18161), 
        .B2(mem_data_out_reg_shift_1[48]), .O(n18201) );
  ND2S U24059 ( .I1(n18359), .I2(mem_data_out_reg_shift_1[64]), .O(n18206) );
  AOI22S U24060 ( .A1(n18165), .A2(mem_data_out_reg_shift_1[40]), .B1(n18357), 
        .B2(mem_data_out_reg_shift_1[88]), .O(n18205) );
  AOI22S U24061 ( .A1(n18168), .A2(mem_data_out_reg_shift_1[8]), .B1(n18169), 
        .B2(mem_data_out_reg_shift_1[96]), .O(n18204) );
  ND3S U24062 ( .I1(n18206), .I2(n18205), .I3(n18204), .O(n18211) );
  ND2S U24063 ( .I1(n18392), .I2(mem_data_out_reg_shift_1[0]), .O(n18209) );
  AOI22S U24064 ( .A1(n18174), .A2(mem_data_out_reg_shift_1[112]), .B1(n18358), 
        .B2(mem_data_out_reg_shift_1[24]), .O(n18208) );
  AOI22S U24065 ( .A1(n18179), .A2(mem_data_out_reg_shift_1[80]), .B1(n18182), 
        .B2(mem_data_out_reg_shift_1[32]), .O(n18207) );
  ND3S U24066 ( .I1(n18209), .I2(n18208), .I3(n18207), .O(n18210) );
  OR3S U24067 ( .I1(n18212), .I2(n18211), .I3(n18210), .O(n15840) );
  AOI22S U24068 ( .A1(n18155), .A2(mem_data_out_reg_shift_1[79]), .B1(n18157), 
        .B2(mem_data_out_reg_shift_1[127]), .O(n18215) );
  AOI22S U24069 ( .A1(n18158), .A2(mem_data_out_reg_shift_1[111]), .B1(n18360), 
        .B2(mem_data_out_reg_shift_1[63]), .O(n18214) );
  AOI22S U24070 ( .A1(n18159), .A2(mem_data_out_reg_shift_1[23]), .B1(n18161), 
        .B2(mem_data_out_reg_shift_1[55]), .O(n18213) );
  ND3S U24071 ( .I1(n18215), .I2(n18214), .I3(n18213), .O(n18224) );
  ND2S U24072 ( .I1(n18359), .I2(mem_data_out_reg_shift_1[71]), .O(n18218) );
  AOI22S U24073 ( .A1(n18165), .A2(mem_data_out_reg_shift_1[47]), .B1(n18357), 
        .B2(mem_data_out_reg_shift_1[95]), .O(n18217) );
  AOI22S U24074 ( .A1(n18168), .A2(mem_data_out_reg_shift_1[15]), .B1(n18169), 
        .B2(mem_data_out_reg_shift_1[103]), .O(n18216) );
  ND2S U24075 ( .I1(n18392), .I2(mem_data_out_reg_shift_1[7]), .O(n18221) );
  AOI22S U24076 ( .A1(n18174), .A2(mem_data_out_reg_shift_1[119]), .B1(n18358), 
        .B2(mem_data_out_reg_shift_1[31]), .O(n18220) );
  AOI22S U24077 ( .A1(n18179), .A2(mem_data_out_reg_shift_1[87]), .B1(n18182), 
        .B2(mem_data_out_reg_shift_1[39]), .O(n18219) );
  ND3S U24078 ( .I1(n18221), .I2(n18220), .I3(n18219), .O(n18222) );
  OR3S U24079 ( .I1(n18224), .I2(n18223), .I3(n18222), .O(n15833) );
  AOI22S U24080 ( .A1(n18155), .A2(mem_data_out_reg_shift_1[75]), .B1(n18157), 
        .B2(mem_data_out_reg_shift_1[123]), .O(n18227) );
  AOI22S U24081 ( .A1(n18158), .A2(mem_data_out_reg_shift_1[107]), .B1(n18360), 
        .B2(mem_data_out_reg_shift_1[59]), .O(n18226) );
  AOI22S U24082 ( .A1(n18159), .A2(mem_data_out_reg_shift_1[19]), .B1(n18161), 
        .B2(mem_data_out_reg_shift_1[51]), .O(n18225) );
  ND3S U24083 ( .I1(n18227), .I2(n18226), .I3(n18225), .O(n18236) );
  ND2S U24084 ( .I1(n18359), .I2(mem_data_out_reg_shift_1[67]), .O(n18230) );
  AOI22S U24085 ( .A1(n18165), .A2(mem_data_out_reg_shift_1[43]), .B1(n18357), 
        .B2(mem_data_out_reg_shift_1[91]), .O(n18229) );
  AOI22S U24086 ( .A1(n18168), .A2(mem_data_out_reg_shift_1[11]), .B1(n18169), 
        .B2(mem_data_out_reg_shift_1[99]), .O(n18228) );
  ND3S U24087 ( .I1(n18230), .I2(n18229), .I3(n18228), .O(n18235) );
  ND2S U24088 ( .I1(n18392), .I2(mem_data_out_reg_shift_1[3]), .O(n18233) );
  AOI22S U24089 ( .A1(n18174), .A2(mem_data_out_reg_shift_1[115]), .B1(n18358), 
        .B2(mem_data_out_reg_shift_1[27]), .O(n18232) );
  AOI22S U24090 ( .A1(n18179), .A2(mem_data_out_reg_shift_1[83]), .B1(n18182), 
        .B2(mem_data_out_reg_shift_1[35]), .O(n18231) );
  ND3S U24091 ( .I1(n18233), .I2(n18232), .I3(n18231), .O(n18234) );
  OR3S U24092 ( .I1(n18236), .I2(n18235), .I3(n18234), .O(n15837) );
  AOI22S U24093 ( .A1(n18155), .A2(mem_data_out_reg_shift_0[76]), .B1(n18157), 
        .B2(mem_data_out_reg_shift_0[124]), .O(n18239) );
  AOI22S U24094 ( .A1(n18158), .A2(mem_data_out_reg_shift_0[108]), .B1(n18360), 
        .B2(mem_data_out_reg_shift_0[60]), .O(n18238) );
  AOI22S U24095 ( .A1(n18159), .A2(mem_data_out_reg_shift_0[20]), .B1(n18161), 
        .B2(mem_data_out_reg_shift_0[52]), .O(n18237) );
  ND3S U24096 ( .I1(n18239), .I2(n18238), .I3(n18237), .O(n18248) );
  ND2S U24097 ( .I1(n18359), .I2(mem_data_out_reg_shift_0[68]), .O(n18242) );
  AOI22S U24098 ( .A1(n18165), .A2(mem_data_out_reg_shift_0[44]), .B1(n18357), 
        .B2(mem_data_out_reg_shift_0[92]), .O(n18241) );
  AOI22S U24099 ( .A1(n18168), .A2(mem_data_out_reg_shift_0[12]), .B1(n18169), 
        .B2(mem_data_out_reg_shift_0[100]), .O(n18240) );
  ND3S U24100 ( .I1(n18242), .I2(n18241), .I3(n18240), .O(n18247) );
  ND2S U24101 ( .I1(n18392), .I2(mem_data_out_reg_shift_0[4]), .O(n18245) );
  AOI22S U24102 ( .A1(n18174), .A2(mem_data_out_reg_shift_0[116]), .B1(n18358), 
        .B2(mem_data_out_reg_shift_0[28]), .O(n18244) );
  AOI22S U24103 ( .A1(n18179), .A2(mem_data_out_reg_shift_0[84]), .B1(n18182), 
        .B2(mem_data_out_reg_shift_0[36]), .O(n18243) );
  ND3S U24104 ( .I1(n18245), .I2(n18244), .I3(n18243), .O(n18246) );
  OR3S U24105 ( .I1(n18248), .I2(n18247), .I3(n18246), .O(n15828) );
  AOI22S U24106 ( .A1(n18155), .A2(mem_data_out_reg_shift_1[76]), .B1(n18157), 
        .B2(mem_data_out_reg_shift_1[124]), .O(n18251) );
  AOI22S U24107 ( .A1(n18158), .A2(mem_data_out_reg_shift_1[108]), .B1(n18360), 
        .B2(mem_data_out_reg_shift_1[60]), .O(n18250) );
  AOI22S U24108 ( .A1(n18159), .A2(mem_data_out_reg_shift_1[20]), .B1(n18161), 
        .B2(mem_data_out_reg_shift_1[52]), .O(n18249) );
  ND2S U24109 ( .I1(n18359), .I2(mem_data_out_reg_shift_1[68]), .O(n18254) );
  AOI22S U24110 ( .A1(n18165), .A2(mem_data_out_reg_shift_1[44]), .B1(n18357), 
        .B2(mem_data_out_reg_shift_1[92]), .O(n18253) );
  AOI22S U24111 ( .A1(n18168), .A2(mem_data_out_reg_shift_1[12]), .B1(n18169), 
        .B2(mem_data_out_reg_shift_1[100]), .O(n18252) );
  ND3S U24112 ( .I1(n18254), .I2(n18253), .I3(n18252), .O(n18259) );
  ND2S U24113 ( .I1(n18392), .I2(mem_data_out_reg_shift_1[4]), .O(n18257) );
  AOI22S U24114 ( .A1(n18174), .A2(mem_data_out_reg_shift_1[116]), .B1(n18358), 
        .B2(mem_data_out_reg_shift_1[28]), .O(n18256) );
  AOI22S U24115 ( .A1(n18179), .A2(mem_data_out_reg_shift_1[84]), .B1(n18182), 
        .B2(mem_data_out_reg_shift_1[36]), .O(n18255) );
  ND3S U24116 ( .I1(n18257), .I2(n18256), .I3(n18255), .O(n18258) );
  OR3S U24117 ( .I1(n18260), .I2(n18259), .I3(n18258), .O(n15836) );
  AOI22S U24118 ( .A1(n18155), .A2(mem_data_out_reg_shift_0[79]), .B1(n18157), 
        .B2(mem_data_out_reg_shift_0[127]), .O(n18263) );
  AOI22S U24119 ( .A1(n18158), .A2(mem_data_out_reg_shift_0[111]), .B1(n18360), 
        .B2(mem_data_out_reg_shift_0[63]), .O(n18262) );
  AOI22S U24120 ( .A1(n18159), .A2(mem_data_out_reg_shift_0[23]), .B1(n18161), 
        .B2(mem_data_out_reg_shift_0[55]), .O(n18261) );
  ND3S U24121 ( .I1(n18263), .I2(n18262), .I3(n18261), .O(n18272) );
  ND2S U24122 ( .I1(n18359), .I2(mem_data_out_reg_shift_0[71]), .O(n18266) );
  AOI22S U24123 ( .A1(n18165), .A2(mem_data_out_reg_shift_0[47]), .B1(n18357), 
        .B2(mem_data_out_reg_shift_0[95]), .O(n18265) );
  AOI22S U24124 ( .A1(n18168), .A2(mem_data_out_reg_shift_0[15]), .B1(n18169), 
        .B2(mem_data_out_reg_shift_0[103]), .O(n18264) );
  ND3S U24125 ( .I1(n18266), .I2(n18265), .I3(n18264), .O(n18271) );
  ND2S U24126 ( .I1(n18392), .I2(mem_data_out_reg_shift_0[7]), .O(n18269) );
  AOI22S U24127 ( .A1(n18174), .A2(mem_data_out_reg_shift_0[119]), .B1(n18358), 
        .B2(mem_data_out_reg_shift_0[31]), .O(n18268) );
  AOI22S U24128 ( .A1(n18179), .A2(mem_data_out_reg_shift_0[87]), .B1(n18182), 
        .B2(mem_data_out_reg_shift_0[39]), .O(n18267) );
  ND3S U24129 ( .I1(n18269), .I2(n18268), .I3(n18267), .O(n18270) );
  OR3S U24130 ( .I1(n18272), .I2(n18271), .I3(n18270), .O(n15825) );
  AOI22S U24131 ( .A1(n18155), .A2(mem_data_out_reg_shift_0[78]), .B1(n18157), 
        .B2(mem_data_out_reg_shift_0[126]), .O(n18275) );
  AOI22S U24132 ( .A1(n18158), .A2(mem_data_out_reg_shift_0[110]), .B1(n18360), 
        .B2(mem_data_out_reg_shift_0[62]), .O(n18274) );
  AOI22S U24133 ( .A1(n18159), .A2(mem_data_out_reg_shift_0[22]), .B1(n18161), 
        .B2(mem_data_out_reg_shift_0[54]), .O(n18273) );
  ND3S U24134 ( .I1(n18275), .I2(n18274), .I3(n18273), .O(n18284) );
  ND2S U24135 ( .I1(n18359), .I2(mem_data_out_reg_shift_0[70]), .O(n18278) );
  AOI22S U24136 ( .A1(n18165), .A2(mem_data_out_reg_shift_0[46]), .B1(n18357), 
        .B2(mem_data_out_reg_shift_0[94]), .O(n18277) );
  AOI22S U24137 ( .A1(n18168), .A2(mem_data_out_reg_shift_0[14]), .B1(n18169), 
        .B2(mem_data_out_reg_shift_0[102]), .O(n18276) );
  ND3S U24138 ( .I1(n18278), .I2(n18277), .I3(n18276), .O(n18283) );
  ND2S U24139 ( .I1(n18392), .I2(mem_data_out_reg_shift_0[6]), .O(n18281) );
  AOI22S U24140 ( .A1(n18174), .A2(mem_data_out_reg_shift_0[118]), .B1(n18358), 
        .B2(mem_data_out_reg_shift_0[30]), .O(n18280) );
  AOI22S U24141 ( .A1(n18179), .A2(mem_data_out_reg_shift_0[86]), .B1(n18182), 
        .B2(mem_data_out_reg_shift_0[38]), .O(n18279) );
  ND3S U24142 ( .I1(n18281), .I2(n18280), .I3(n18279), .O(n18282) );
  OR3S U24143 ( .I1(n18284), .I2(n18283), .I3(n18282), .O(n15826) );
  AOI22S U24144 ( .A1(n18155), .A2(mem_data_out_reg_shift_1[73]), .B1(n18157), 
        .B2(mem_data_out_reg_shift_1[121]), .O(n18287) );
  AOI22S U24145 ( .A1(n18158), .A2(mem_data_out_reg_shift_1[105]), .B1(n18360), 
        .B2(mem_data_out_reg_shift_1[57]), .O(n18286) );
  AOI22S U24146 ( .A1(n18159), .A2(mem_data_out_reg_shift_1[17]), .B1(n18161), 
        .B2(mem_data_out_reg_shift_1[49]), .O(n18285) );
  ND3S U24147 ( .I1(n18287), .I2(n18286), .I3(n18285), .O(n18296) );
  ND2S U24148 ( .I1(n18359), .I2(mem_data_out_reg_shift_1[65]), .O(n18290) );
  AOI22S U24149 ( .A1(n18165), .A2(mem_data_out_reg_shift_1[41]), .B1(n18357), 
        .B2(mem_data_out_reg_shift_1[89]), .O(n18289) );
  AOI22S U24150 ( .A1(n18168), .A2(mem_data_out_reg_shift_1[9]), .B1(n18169), 
        .B2(mem_data_out_reg_shift_1[97]), .O(n18288) );
  ND3S U24151 ( .I1(n18290), .I2(n18289), .I3(n18288), .O(n18295) );
  ND2S U24152 ( .I1(n18392), .I2(mem_data_out_reg_shift_1[1]), .O(n18293) );
  AOI22S U24153 ( .A1(n18174), .A2(mem_data_out_reg_shift_1[113]), .B1(n18358), 
        .B2(mem_data_out_reg_shift_1[25]), .O(n18292) );
  AOI22S U24154 ( .A1(n18179), .A2(mem_data_out_reg_shift_1[81]), .B1(n18182), 
        .B2(mem_data_out_reg_shift_1[33]), .O(n18291) );
  OR3S U24155 ( .I1(n18296), .I2(n18295), .I3(n18294), .O(n15839) );
  AOI22S U24156 ( .A1(n18155), .A2(mem_data_out_reg_shift_0[77]), .B1(n18157), 
        .B2(mem_data_out_reg_shift_0[125]), .O(n18299) );
  AOI22S U24157 ( .A1(n18158), .A2(mem_data_out_reg_shift_0[109]), .B1(n18360), 
        .B2(mem_data_out_reg_shift_0[61]), .O(n18298) );
  AOI22S U24158 ( .A1(n18159), .A2(mem_data_out_reg_shift_0[21]), .B1(n18161), 
        .B2(mem_data_out_reg_shift_0[53]), .O(n18297) );
  ND3S U24159 ( .I1(n18299), .I2(n18298), .I3(n18297), .O(n18308) );
  ND2S U24160 ( .I1(n18359), .I2(mem_data_out_reg_shift_0[69]), .O(n18302) );
  AOI22S U24161 ( .A1(n18165), .A2(mem_data_out_reg_shift_0[45]), .B1(n18357), 
        .B2(mem_data_out_reg_shift_0[93]), .O(n18301) );
  AOI22S U24162 ( .A1(n18168), .A2(mem_data_out_reg_shift_0[13]), .B1(n18169), 
        .B2(mem_data_out_reg_shift_0[101]), .O(n18300) );
  ND3S U24163 ( .I1(n18302), .I2(n18301), .I3(n18300), .O(n18307) );
  ND2S U24164 ( .I1(n18392), .I2(mem_data_out_reg_shift_0[5]), .O(n18305) );
  AOI22S U24165 ( .A1(n18174), .A2(mem_data_out_reg_shift_0[117]), .B1(n18358), 
        .B2(mem_data_out_reg_shift_0[29]), .O(n18304) );
  AOI22S U24166 ( .A1(n18179), .A2(mem_data_out_reg_shift_0[85]), .B1(n18182), 
        .B2(mem_data_out_reg_shift_0[37]), .O(n18303) );
  ND3S U24167 ( .I1(n18305), .I2(n18304), .I3(n18303), .O(n18306) );
  OR3S U24168 ( .I1(n18308), .I2(n18307), .I3(n18306), .O(n15827) );
  AOI22S U24169 ( .A1(n18155), .A2(mem_data_out_reg_shift_0[72]), .B1(n18157), 
        .B2(mem_data_out_reg_shift_0[120]), .O(n18311) );
  AOI22S U24170 ( .A1(n18158), .A2(mem_data_out_reg_shift_0[104]), .B1(n18360), 
        .B2(mem_data_out_reg_shift_0[56]), .O(n18310) );
  AOI22S U24171 ( .A1(n18159), .A2(mem_data_out_reg_shift_0[16]), .B1(n18161), 
        .B2(mem_data_out_reg_shift_0[48]), .O(n18309) );
  ND3S U24172 ( .I1(n18311), .I2(n18310), .I3(n18309), .O(n18320) );
  ND2S U24173 ( .I1(n18359), .I2(mem_data_out_reg_shift_0[64]), .O(n18314) );
  AOI22S U24174 ( .A1(n18165), .A2(mem_data_out_reg_shift_0[40]), .B1(n18357), 
        .B2(mem_data_out_reg_shift_0[88]), .O(n18313) );
  AOI22S U24175 ( .A1(n18168), .A2(mem_data_out_reg_shift_0[8]), .B1(n18169), 
        .B2(mem_data_out_reg_shift_0[96]), .O(n18312) );
  ND3S U24176 ( .I1(n18314), .I2(n18313), .I3(n18312), .O(n18319) );
  ND2S U24177 ( .I1(n18392), .I2(mem_data_out_reg_shift_0[0]), .O(n18317) );
  AOI22S U24178 ( .A1(n18174), .A2(mem_data_out_reg_shift_0[112]), .B1(n18358), 
        .B2(mem_data_out_reg_shift_0[24]), .O(n18316) );
  AOI22S U24179 ( .A1(n18179), .A2(mem_data_out_reg_shift_0[80]), .B1(n18182), 
        .B2(mem_data_out_reg_shift_0[32]), .O(n18315) );
  ND3S U24180 ( .I1(n18317), .I2(n18316), .I3(n18315), .O(n18318) );
  OR3S U24181 ( .I1(n18320), .I2(n18319), .I3(n18318), .O(n15832) );
  AOI22S U24182 ( .A1(n18155), .A2(mem_data_out_reg_shift_1[78]), .B1(n18157), 
        .B2(mem_data_out_reg_shift_1[126]), .O(n18323) );
  AOI22S U24183 ( .A1(n18158), .A2(mem_data_out_reg_shift_1[110]), .B1(n18360), 
        .B2(mem_data_out_reg_shift_1[62]), .O(n18322) );
  AOI22S U24184 ( .A1(n18159), .A2(mem_data_out_reg_shift_1[22]), .B1(n18161), 
        .B2(mem_data_out_reg_shift_1[54]), .O(n18321) );
  ND3S U24185 ( .I1(n18323), .I2(n18322), .I3(n18321), .O(n18332) );
  ND2S U24186 ( .I1(n18359), .I2(mem_data_out_reg_shift_1[70]), .O(n18326) );
  AOI22S U24187 ( .A1(n18165), .A2(mem_data_out_reg_shift_1[46]), .B1(n18357), 
        .B2(mem_data_out_reg_shift_1[94]), .O(n18325) );
  AOI22S U24188 ( .A1(n18168), .A2(mem_data_out_reg_shift_1[14]), .B1(n18169), 
        .B2(mem_data_out_reg_shift_1[102]), .O(n18324) );
  ND3S U24189 ( .I1(n18326), .I2(n18325), .I3(n18324), .O(n18331) );
  ND2S U24190 ( .I1(n18392), .I2(mem_data_out_reg_shift_1[6]), .O(n18329) );
  AOI22S U24191 ( .A1(n18174), .A2(mem_data_out_reg_shift_1[118]), .B1(n18358), 
        .B2(mem_data_out_reg_shift_1[30]), .O(n18328) );
  AOI22S U24192 ( .A1(n18179), .A2(mem_data_out_reg_shift_1[86]), .B1(n18182), 
        .B2(mem_data_out_reg_shift_1[38]), .O(n18327) );
  ND3S U24193 ( .I1(n18329), .I2(n18328), .I3(n18327), .O(n18330) );
  OR3S U24194 ( .I1(n18332), .I2(n18331), .I3(n18330), .O(n15834) );
  AOI22S U24195 ( .A1(n18155), .A2(mem_data_out_reg_shift_1[74]), .B1(n18157), 
        .B2(mem_data_out_reg_shift_1[122]), .O(n18335) );
  AOI22S U24196 ( .A1(n18158), .A2(mem_data_out_reg_shift_1[106]), .B1(n18360), 
        .B2(mem_data_out_reg_shift_1[58]), .O(n18334) );
  AOI22S U24197 ( .A1(n18159), .A2(mem_data_out_reg_shift_1[18]), .B1(n18161), 
        .B2(mem_data_out_reg_shift_1[50]), .O(n18333) );
  ND3S U24198 ( .I1(n18335), .I2(n18334), .I3(n18333), .O(n18344) );
  ND2S U24199 ( .I1(n18359), .I2(mem_data_out_reg_shift_1[66]), .O(n18338) );
  AOI22S U24200 ( .A1(n18165), .A2(mem_data_out_reg_shift_1[42]), .B1(n18357), 
        .B2(mem_data_out_reg_shift_1[90]), .O(n18337) );
  AOI22S U24201 ( .A1(n18168), .A2(mem_data_out_reg_shift_1[10]), .B1(n18169), 
        .B2(mem_data_out_reg_shift_1[98]), .O(n18336) );
  ND3S U24202 ( .I1(n18338), .I2(n18337), .I3(n18336), .O(n18343) );
  ND2S U24203 ( .I1(n18392), .I2(mem_data_out_reg_shift_1[2]), .O(n18341) );
  AOI22S U24204 ( .A1(n18174), .A2(mem_data_out_reg_shift_1[114]), .B1(n18358), 
        .B2(mem_data_out_reg_shift_1[26]), .O(n18340) );
  AOI22S U24205 ( .A1(n18179), .A2(mem_data_out_reg_shift_1[82]), .B1(n18182), 
        .B2(mem_data_out_reg_shift_1[34]), .O(n18339) );
  ND3S U24206 ( .I1(n18341), .I2(n18340), .I3(n18339), .O(n18342) );
  OR3S U24207 ( .I1(n18344), .I2(n18343), .I3(n18342), .O(n15838) );
  AOI22S U24208 ( .A1(n18155), .A2(mem_data_out_reg_shift_1[77]), .B1(n18157), 
        .B2(mem_data_out_reg_shift_1[125]), .O(n18347) );
  AOI22S U24209 ( .A1(n18158), .A2(mem_data_out_reg_shift_1[109]), .B1(n18360), 
        .B2(mem_data_out_reg_shift_1[61]), .O(n18346) );
  AOI22S U24210 ( .A1(n18159), .A2(mem_data_out_reg_shift_1[21]), .B1(n18161), 
        .B2(mem_data_out_reg_shift_1[53]), .O(n18345) );
  ND3S U24211 ( .I1(n18347), .I2(n18346), .I3(n18345), .O(n18356) );
  ND2S U24212 ( .I1(n18359), .I2(mem_data_out_reg_shift_1[69]), .O(n18350) );
  AOI22S U24213 ( .A1(n18165), .A2(mem_data_out_reg_shift_1[45]), .B1(n18357), 
        .B2(mem_data_out_reg_shift_1[93]), .O(n18349) );
  AOI22S U24214 ( .A1(n18168), .A2(mem_data_out_reg_shift_1[13]), .B1(n18169), 
        .B2(mem_data_out_reg_shift_1[101]), .O(n18348) );
  ND3S U24215 ( .I1(n18350), .I2(n18349), .I3(n18348), .O(n18355) );
  ND2S U24216 ( .I1(n18392), .I2(mem_data_out_reg_shift_1[5]), .O(n18353) );
  AOI22S U24217 ( .A1(n18174), .A2(mem_data_out_reg_shift_1[117]), .B1(n18358), 
        .B2(mem_data_out_reg_shift_1[29]), .O(n18352) );
  AOI22S U24218 ( .A1(n18179), .A2(mem_data_out_reg_shift_1[85]), .B1(n18182), 
        .B2(mem_data_out_reg_shift_1[37]), .O(n18351) );
  ND3S U24219 ( .I1(n18353), .I2(n18352), .I3(n18351), .O(n18354) );
  OR3S U24220 ( .I1(n18356), .I2(n18355), .I3(n18354), .O(n15835) );
  AOI22S U24221 ( .A1(n18157), .A2(mem_data_out_reg_shift_0[121]), .B1(n18357), 
        .B2(mem_data_out_reg_shift_0[89]), .O(n18371) );
  AOI22S U24222 ( .A1(n18155), .A2(mem_data_out_reg_shift_0[73]), .B1(n18165), 
        .B2(mem_data_out_reg_shift_0[41]), .O(n18370) );
  AOI22S U24223 ( .A1(n18159), .A2(mem_data_out_reg_shift_0[17]), .B1(n18358), 
        .B2(mem_data_out_reg_shift_0[25]), .O(n18368) );
  AOI22S U24224 ( .A1(n18179), .A2(mem_data_out_reg_shift_0[81]), .B1(n18182), 
        .B2(mem_data_out_reg_shift_0[33]), .O(n18367) );
  ND2S U24225 ( .I1(n18359), .I2(mem_data_out_reg_shift_0[65]), .O(n18366) );
  AOI22S U24226 ( .A1(n18161), .A2(mem_data_out_reg_shift_0[49]), .B1(n18360), 
        .B2(mem_data_out_reg_shift_0[57]), .O(n18363) );
  AOI22S U24227 ( .A1(n18174), .A2(mem_data_out_reg_shift_0[113]), .B1(n18158), 
        .B2(mem_data_out_reg_shift_0[105]), .O(n18362) );
  AOI22S U24228 ( .A1(n18168), .A2(mem_data_out_reg_shift_0[9]), .B1(n18169), 
        .B2(mem_data_out_reg_shift_0[97]), .O(n18361) );
  ND3S U24229 ( .I1(n18363), .I2(n18362), .I3(n18361), .O(n18364) );
  AO12S U24230 ( .B1(n18392), .B2(mem_data_out_reg_shift_0[1]), .A1(n18364), 
        .O(n18365) );
  AN4B1S U24231 ( .I1(n18368), .I2(n18367), .I3(n18366), .B1(n18365), .O(
        n18369) );
  ND3S U24232 ( .I1(n18371), .I2(n18370), .I3(n18369), .O(n15831) );
  NR2 U24233 ( .I1(medfilt_state[1]), .I2(medfilt_state[2]), .O(n18373) );
  NR2 U24234 ( .I1(cnt_bdyn[1]), .I2(n30372), .O(n30132) );
  INV1S U24235 ( .I(cnt_bdyn[2]), .O(n30365) );
  NR2 U24236 ( .I1(n21156), .I2(n21138), .O(n22769) );
  INV1S U24237 ( .I(cnt_dyn[3]), .O(n30307) );
  ND2S U24238 ( .I1(n30305), .I2(n30307), .O(n30281) );
  NR2 U24239 ( .I1(cnt_bdyn[5]), .I2(cnt_bdyn[4]), .O(n30321) );
  INV1S U24240 ( .I(cnt_bdyn[7]), .O(n30353) );
  INV1S U24241 ( .I(cnt_bdyn[6]), .O(n30323) );
  NR2 U24242 ( .I1(n30281), .I2(n30129), .O(n18463) );
  INV1S U24243 ( .I(cnt_bdyn[8]), .O(n30280) );
  INV3 U24244 ( .I(medfilt_state[0]), .O(n19088) );
  AO13S U24245 ( .B1(n15918), .B2(n18463), .B3(n30280), .A1(n19088), .O(n18372) );
  NR2 U24246 ( .I1(medfilt_state[3]), .I2(n30360), .O(n24925) );
  AO13S U24247 ( .B1(n24942), .B2(n18373), .B3(n18372), .A1(n24925), .O(n19091) );
  INV2 U24248 ( .I(medfilt_state[3]), .O(n30242) );
  ND3P U24249 ( .I1(n18373), .I2(n30242), .I3(n19088), .O(n23993) );
  BUF6 U24250 ( .I(n23993), .O(n24047) );
  INV3 U24251 ( .I(medfilt_state[2]), .O(n18374) );
  NR2F U24252 ( .I1(medfilt_state[1]), .I2(n18374), .O(n24928) );
  ND2 U24253 ( .I1(n24928), .I2(n19088), .O(n24068) );
  OR2 U24254 ( .I1(medfilt_state[2]), .I2(n19088), .O(n23685) );
  NR2P U24255 ( .I1(n30453), .I2(n23685), .O(n24909) );
  INV1S U24256 ( .I(n24909), .O(n24923) );
  NR2 U24257 ( .I1(n18385), .I2(n18375), .O(n18386) );
  XOR2HS U24258 ( .I1(medfilt_cnt[1]), .I2(n18386), .O(n18377) );
  ND2S U24259 ( .I1(n18383), .I2(medfilt_cnt[3]), .O(n18376) );
  ND2S U24260 ( .I1(n18377), .I2(n18376), .O(n18378) );
  NR2 U24261 ( .I1(n18392), .I2(n18378), .O(n18382) );
  INV1S U24262 ( .I(medfilt_cnt[2]), .O(n30246) );
  XNR2HS U24263 ( .I1(cnt_dyn_base[2]), .I2(n30246), .O(n24907) );
  XNR2HS U24264 ( .I1(n18385), .I2(n24907), .O(n18381) );
  XNR2HS U24265 ( .I1(cnt_dyn_base[0]), .I2(medfilt_cnt[0]), .O(n24906) );
  XNR2HS U24266 ( .I1(cnt_dyn_base[3]), .I2(medfilt_cnt[3]), .O(n24905) );
  NR2 U24267 ( .I1(n24905), .I2(n18383), .O(n18379) );
  NR2 U24268 ( .I1(n24906), .I2(n18379), .O(n18380) );
  ND3S U24269 ( .I1(n18382), .I2(n18381), .I3(n18380), .O(n24922) );
  MUX2S U24270 ( .A(n24068), .B(n24923), .S(n24922), .O(n18395) );
  NR2 U24271 ( .I1(n19088), .I2(n24922), .O(n19089) );
  OR2S U24272 ( .I1(n24919), .I2(n19089), .O(n24932) );
  NR2 U24273 ( .I1(n24903), .I2(n18383), .O(n18384) );
  XOR2HS U24274 ( .I1(medfilt_cnt2[3]), .I2(n18384), .O(n18391) );
  XNR3S U24275 ( .I1(cnt_dyn_base[2]), .I2(medfilt_cnt2[2]), .I3(n18385), .O(
        n18389) );
  XOR2HS U24276 ( .I1(medfilt_cnt2[1]), .I2(n18386), .O(n18388) );
  INV1S U24277 ( .I(medfilt_cnt2[0]), .O(n30427) );
  XNR2HS U24278 ( .I1(n30427), .I2(cnt_dyn_base[0]), .O(n18387) );
  ND3S U24279 ( .I1(n18389), .I2(n18388), .I3(n18387), .O(n18390) );
  NR3 U24280 ( .I1(n18392), .I2(n18391), .I3(n18390), .O(n24929) );
  INV1 U24281 ( .I(medfilt_state[1]), .O(n23637) );
  ND2S U24282 ( .I1(n24929), .I2(n24118), .O(n18393) );
  ND2S U24283 ( .I1(n24928), .I2(medfilt_state[0]), .O(n23684) );
  ND2T U24284 ( .I1(n24118), .I2(n23684), .O(n30241) );
  ND2S U24285 ( .I1(n18393), .I2(n30241), .O(n18394) );
  AO13S U24286 ( .B1(n18395), .B2(n24932), .B3(n18394), .A1(medfilt_state[3]), 
        .O(n18396) );
  NR2 U24287 ( .I1(cs[1]), .I2(n18397), .O(n24934) );
  INV1S U24288 ( .I(n24934), .O(n24936) );
  ND2S U24289 ( .I1(n24936), .I2(n24897), .O(n30412) );
  INV1S U24290 ( .I(n30412), .O(n18399) );
  ND2S U24291 ( .I1(n18399), .I2(n18398), .O(n15789) );
  ND2S U24292 ( .I1(action_reg[16]), .I2(n18401), .O(n18405) );
  OR3S U24293 ( .I1(cnt[7]), .I2(cnt[6]), .I3(cnt[4]), .O(n18402) );
  NR3 U24294 ( .I1(cnt[3]), .I2(cnt[5]), .I3(n18402), .O(n30429) );
  ND2S U24295 ( .I1(n30429), .I2(n24967), .O(n18403) );
  NR2 U24296 ( .I1(n24934), .I2(n18401), .O(n18418) );
  INV1S U24297 ( .I(cnt[2]), .O(n30259) );
  OA12S U24298 ( .B1(cnt[1]), .B2(n30259), .A1(n18418), .O(n18426) );
  NR2 U24299 ( .I1(n30400), .I2(n18426), .O(n18408) );
  ND2S U24300 ( .I1(n24967), .I2(action_in_reg[1]), .O(n30403) );
  MOAI1S U24301 ( .A1(n18408), .A2(action_reg[13]), .B1(n18408), .B2(n30403), 
        .O(n18404) );
  ND2S U24302 ( .I1(n18405), .I2(n18404), .O(n15777) );
  ND2S U24303 ( .I1(action_reg[17]), .I2(n18401), .O(n18407) );
  ND2S U24304 ( .I1(n24967), .I2(action_in_reg[2]), .O(n30406) );
  MOAI1S U24305 ( .A1(n18408), .A2(action_reg[14]), .B1(n18408), .B2(n30406), 
        .O(n18406) );
  ND2S U24306 ( .I1(n18407), .I2(n18406), .O(n15769) );
  ND2S U24307 ( .I1(action_reg[15]), .I2(n18401), .O(n18410) );
  ND2S U24308 ( .I1(n24967), .I2(action_in_reg[0]), .O(n30401) );
  MOAI1S U24309 ( .A1(n18408), .A2(action_reg[12]), .B1(n18408), .B2(n30401), 
        .O(n18409) );
  ND2S U24310 ( .I1(n18410), .I2(n18409), .O(n15785) );
  ND2S U24311 ( .I1(action_reg[3]), .I2(n18401), .O(n18412) );
  OA12S U24312 ( .B1(cnt[1]), .B2(cnt[2]), .A1(n18418), .O(n18434) );
  NR2 U24313 ( .I1(n30400), .I2(n18434), .O(n18415) );
  MOAI1S U24314 ( .A1(n18415), .A2(action_reg[0]), .B1(n18415), .B2(n30401), 
        .O(n18411) );
  ND2S U24315 ( .I1(n18412), .I2(n18411), .O(n15781) );
  ND2S U24316 ( .I1(action_reg[4]), .I2(n18401), .O(n18414) );
  MOAI1S U24317 ( .A1(n18415), .A2(action_reg[1]), .B1(n18415), .B2(n30403), 
        .O(n18413) );
  ND2S U24318 ( .I1(n18414), .I2(n18413), .O(n15773) );
  ND2S U24319 ( .I1(action_reg[5]), .I2(n18401), .O(n18417) );
  MOAI1S U24320 ( .A1(n18415), .A2(action_reg[2]), .B1(n18415), .B2(n30406), 
        .O(n18416) );
  ND2S U24321 ( .I1(n18417), .I2(n18416), .O(n15765) );
  ND2S U24322 ( .I1(action_reg[10]), .I2(n18401), .O(n18420) );
  INV1S U24323 ( .I(n18418), .O(n30397) );
  OAI22S U24324 ( .A1(cnt[1]), .A2(n30397), .B1(n30259), .B2(n30397), .O(
        n18429) );
  NR2 U24325 ( .I1(n30400), .I2(n18429), .O(n18423) );
  MOAI1S U24326 ( .A1(n18423), .A2(action_reg[7]), .B1(n18423), .B2(n30403), 
        .O(n18419) );
  ND2S U24327 ( .I1(n18420), .I2(n18419), .O(n15775) );
  ND2S U24328 ( .I1(action_reg[11]), .I2(n18401), .O(n18422) );
  MOAI1S U24329 ( .A1(n18423), .A2(action_reg[8]), .B1(n18423), .B2(n30406), 
        .O(n18421) );
  ND2S U24330 ( .I1(n18422), .I2(n18421), .O(n15767) );
  ND2S U24331 ( .I1(action_reg[9]), .I2(n18401), .O(n18425) );
  MOAI1S U24332 ( .A1(n18423), .A2(action_reg[6]), .B1(n18423), .B2(n30401), 
        .O(n18424) );
  ND2S U24333 ( .I1(n18425), .I2(n18424), .O(n15783) );
  ND2S U24334 ( .I1(action_reg[18]), .I2(n18401), .O(n18428) );
  AOI13HS U24335 ( .B1(cnt[0]), .B2(n30429), .B3(n24967), .A1(n30397), .O(
        n30398) );
  NR2 U24336 ( .I1(n30398), .I2(n18426), .O(n18441) );
  MOAI1S U24337 ( .A1(n18441), .A2(action_reg[15]), .B1(n18441), .B2(n30401), 
        .O(n18427) );
  ND2S U24338 ( .I1(n18428), .I2(n18427), .O(n15786) );
  ND2S U24339 ( .I1(action_reg[13]), .I2(n18401), .O(n18431) );
  NR2 U24340 ( .I1(n30398), .I2(n18429), .O(n18444) );
  MOAI1S U24341 ( .A1(n18444), .A2(action_reg[10]), .B1(n18444), .B2(n30403), 
        .O(n18430) );
  ND2S U24342 ( .I1(n18431), .I2(n18430), .O(n15776) );
  ND2S U24343 ( .I1(action_reg[14]), .I2(n18401), .O(n18433) );
  MOAI1S U24344 ( .A1(n18444), .A2(action_reg[11]), .B1(n18444), .B2(n30406), 
        .O(n18432) );
  ND2S U24345 ( .I1(n18433), .I2(n18432), .O(n15768) );
  ND2S U24346 ( .I1(action_reg[8]), .I2(n18401), .O(n18436) );
  NR2 U24347 ( .I1(n30398), .I2(n18434), .O(n18447) );
  MOAI1S U24348 ( .A1(n18447), .A2(action_reg[5]), .B1(n18447), .B2(n30406), 
        .O(n18435) );
  ND2S U24349 ( .I1(n18436), .I2(n18435), .O(n15766) );
  ND2S U24350 ( .I1(action_reg[6]), .I2(n18401), .O(n18438) );
  MOAI1S U24351 ( .A1(n18447), .A2(action_reg[3]), .B1(n18447), .B2(n30401), 
        .O(n18437) );
  ND2S U24352 ( .I1(n18438), .I2(n18437), .O(n15782) );
  ND2S U24353 ( .I1(action_reg[20]), .I2(n18401), .O(n18440) );
  MOAI1S U24354 ( .A1(n18441), .A2(action_reg[17]), .B1(n18441), .B2(n30406), 
        .O(n18439) );
  ND2S U24355 ( .I1(n18440), .I2(n18439), .O(n15770) );
  ND2S U24356 ( .I1(action_reg[19]), .I2(n18401), .O(n18443) );
  MOAI1S U24357 ( .A1(n18441), .A2(action_reg[16]), .B1(n18441), .B2(n30403), 
        .O(n18442) );
  ND2S U24358 ( .I1(n18443), .I2(n18442), .O(n15778) );
  ND2S U24359 ( .I1(action_reg[12]), .I2(n18401), .O(n18446) );
  MOAI1S U24360 ( .A1(n18444), .A2(action_reg[9]), .B1(n18444), .B2(n30401), 
        .O(n18445) );
  ND2S U24361 ( .I1(n18446), .I2(n18445), .O(n15784) );
  ND2S U24362 ( .I1(action_reg[7]), .I2(n18401), .O(n18449) );
  MOAI1S U24363 ( .A1(n18447), .A2(action_reg[4]), .B1(n18447), .B2(n30403), 
        .O(n18448) );
  ND2S U24364 ( .I1(n18449), .I2(n18448), .O(n15774) );
  NR2 U24365 ( .I1(cnt_bdyn[1]), .I2(cnt_bdyn[0]), .O(n30303) );
  NR2 U24366 ( .I1(n30306), .I2(cnt_bdyn[3]), .O(n30322) );
  NR2 U24367 ( .I1(cnt_dyn[1]), .I2(cnt_dyn[0]), .O(n30299) );
  AN2 U24368 ( .I1(n30322), .I2(n30299), .O(n22893) );
  ND2S U24369 ( .I1(n18450), .I2(n29427), .O(n18462) );
  INV1S U24370 ( .I(cnt_dyn[0]), .O(n30333) );
  XOR2HS U24371 ( .I1(cnt_dyn_base[2]), .I2(n30365), .O(n18451) );
  OA12S U24372 ( .B1(n30333), .B2(cnt_bdyn[0]), .A1(n18451), .O(n18454) );
  MUX2S U24373 ( .A(cnt_dyn[0]), .B(n30372), .S(n24898), .O(n18452) );
  ND3S U24374 ( .I1(n18454), .I2(n18453), .I3(n18452), .O(n18460) );
  XOR2HS U24375 ( .I1(cnt_dyn_base[3]), .I2(n30330), .O(n18457) );
  XOR2HS U24376 ( .I1(cnt_dyn_base[1]), .I2(n30369), .O(n18456) );
  ND3S U24377 ( .I1(n18642), .I2(n18457), .I3(n18456), .O(n18459) );
  AN2B1S U24378 ( .I1(out_valid), .B1(out_valid_a1), .O(n30432) );
  NR2 U24379 ( .I1(n30409), .I2(n18458), .O(n30379) );
  MOAI1S U24380 ( .A1(n18460), .A2(n18459), .B1(n30432), .B2(n30379), .O(
        n18461) );
  AOI13HS U24381 ( .B1(n22893), .B2(n18463), .B3(n18462), .A1(n18461), .O(
        n18466) );
  BUF2 U24382 ( .I(n18464), .O(n24100) );
  ND3S U24383 ( .I1(n19127), .I2(n24100), .I3(medfilt_state[3]), .O(n18465) );
  ND2S U24384 ( .I1(n18466), .I2(n18465), .O(n15795) );
  AOI22S U24385 ( .A1(action_done), .A2(n30383), .B1(in_valid), .B2(n24934), 
        .O(n18468) );
  INV1S U24386 ( .I(in_valid2), .O(n30257) );
  NR2 U24387 ( .I1(in_valid2), .I2(n30390), .O(n30389) );
  AOI13HS U24388 ( .B1(last_in_valid2), .B2(n24967), .B3(n30257), .A1(n30389), 
        .O(n18467) );
  ND2S U24389 ( .I1(n18468), .I2(n18467), .O(n15793) );
  ND2S U24390 ( .I1(cnt_20[0]), .I2(cnt_20[1]), .O(n30227) );
  OA112S U24391 ( .C1(cnt_20[0]), .C2(cnt_20[1]), .A1(n24942), .B1(n30227), 
        .O(cnt_20_n[1]) );
  INV1S U24392 ( .I(n25194), .O(n20322) );
  NR2 U24393 ( .I1(n18579), .I2(n18567), .O(n25065) );
  MOAI1S U24394 ( .A1(n20322), .A2(n25066), .B1(n25193), .B2(n25065), .O(
        n18471) );
  MUX2S U24395 ( .A(n30005), .B(n20156), .S(gray_img[1827]), .O(n18473) );
  ND2S U24396 ( .I1(n18473), .I2(n18472), .O(n14705) );
  INV1S U24397 ( .I(medfilt_out_reg[1]), .O(n18474) );
  NR2 U24398 ( .I1(n18474), .I2(n18734), .O(n18475) );
  AN2B1S U24399 ( .I1(medfilt_cnt_d1[3]), .B1(n18476), .O(n18641) );
  NR2 U24400 ( .I1(n18820), .I2(n25049), .O(n19720) );
  INV1S U24401 ( .I(n19720), .O(n18829) );
  NR2 U24402 ( .I1(n18533), .I2(n18578), .O(n25057) );
  MOAI1S U24403 ( .A1(n18829), .A2(n25058), .B1(n19719), .B2(n25057), .O(
        n18479) );
  INV2 U24404 ( .I(n27447), .O(n29597) );
  ND2S U24405 ( .I1(n18481), .I2(n18480), .O(n14310) );
  INV1S U24406 ( .I(medfilt_out_reg[2]), .O(n18482) );
  NR2 U24407 ( .I1(n18482), .I2(n18734), .O(n18483) );
  NR2 U24408 ( .I1(n18542), .I2(n18571), .O(n25162) );
  INV1S U24409 ( .I(n25162), .O(n25362) );
  NR2 U24410 ( .I1(n18543), .I2(n18572), .O(n25361) );
  MOAI1S U24411 ( .A1(n25362), .A2(n18829), .B1(n25361), .B2(n19719), .O(
        n18484) );
  INV2 U24412 ( .I(n27447), .O(n30050) );
  ND2S U24413 ( .I1(n18486), .I2(n18485), .O(n14647) );
  INV1S U24414 ( .I(n25372), .O(n25367) );
  MOAI1S U24415 ( .A1(n25367), .A2(n18829), .B1(n25370), .B2(n19719), .O(
        n18487) );
  ND2S U24416 ( .I1(n18489), .I2(n18488), .O(n14639) );
  INV2 U24417 ( .I(n27447), .O(n29587) );
  ND2S U24418 ( .I1(n18491), .I2(n18490), .O(n14711) );
  NR2 U24419 ( .I1(n18533), .I2(n18567), .O(n25053) );
  MOAI1S U24420 ( .A1(n18829), .A2(n25054), .B1(n19719), .B2(n25053), .O(
        n18492) );
  ND2S U24421 ( .I1(n18494), .I2(n18493), .O(n14727) );
  MOAI1S U24422 ( .A1(n18829), .A2(n25066), .B1(n19719), .B2(n25065), .O(
        n18495) );
  INV2 U24423 ( .I(n27447), .O(n29566) );
  ND2S U24424 ( .I1(n18497), .I2(n18496), .O(n14695) );
  INV2 U24425 ( .I(n27447), .O(n30044) );
  ND2S U24426 ( .I1(n18499), .I2(n18498), .O(n14446) );
  ND2S U24427 ( .I1(n18501), .I2(n18500), .O(n14326) );
  ND2S U24428 ( .I1(n18503), .I2(n18502), .O(n14294) );
  NR2 U24429 ( .I1(n18509), .I2(n18576), .O(n19758) );
  INV1S U24430 ( .I(n19758), .O(n25297) );
  NR2 U24431 ( .I1(n18510), .I2(n18578), .O(n25296) );
  MOAI1S U24432 ( .A1(n20322), .A2(n25297), .B1(n25193), .B2(n25296), .O(
        n18504) );
  ND2S U24433 ( .I1(n18506), .I2(n18505), .O(n14785) );
  ND2S U24434 ( .I1(n18508), .I2(n18507), .O(n14384) );
  NR2 U24435 ( .I1(n18509), .I2(n18566), .O(n19772) );
  INV1S U24436 ( .I(n19772), .O(n25301) );
  NR2 U24437 ( .I1(n18510), .I2(n18567), .O(n25300) );
  MOAI1S U24438 ( .A1(n20322), .A2(n25301), .B1(n25193), .B2(n25300), .O(
        n18511) );
  ND2S U24439 ( .I1(n18513), .I2(n18512), .O(n14400) );
  ND2S U24440 ( .I1(n18515), .I2(n18514), .O(n14801) );
  INV2 U24441 ( .I(n27447), .O(n30056) );
  MOAI1S U24442 ( .A1(n20322), .A2(n25058), .B1(n25193), .B2(n25057), .O(
        n18516) );
  INV1S U24443 ( .I(medfilt_out_reg[5]), .O(n18517) );
  NR2 U24444 ( .I1(n18517), .I2(n18734), .O(n18518) );
  ND2S U24445 ( .I1(n15891), .I2(n20787), .O(n18519) );
  ND2S U24446 ( .I1(n18520), .I2(n18519), .O(n15120) );
  MOAI1S U24447 ( .A1(n20322), .A2(n25054), .B1(n25193), .B2(n25053), .O(
        n18521) );
  ND2S U24448 ( .I1(n15891), .I2(n20824), .O(n18522) );
  ND2S U24449 ( .I1(n18523), .I2(n18522), .O(n15136) );
  ND2S U24450 ( .I1(n27751), .I2(n20522), .O(n18525) );
  ND2S U24451 ( .I1(n18525), .I2(n18524), .O(n15246) );
  ND2S U24452 ( .I1(n15891), .I2(n20541), .O(n18527) );
  MUX2S U24453 ( .A(n29032), .B(n20541), .S(gray_img[1781]), .O(n18526) );
  ND2S U24454 ( .I1(n18527), .I2(n18526), .O(n15110) );
  INV1S U24455 ( .I(n29831), .O(n27751) );
  ND2S U24456 ( .I1(n27751), .I2(n20477), .O(n18529) );
  ND2S U24457 ( .I1(n18529), .I2(n18528), .O(n15238) );
  ND2S U24458 ( .I1(n15891), .I2(n20063), .O(n18531) );
  ND2S U24459 ( .I1(n18531), .I2(n18530), .O(n15094) );
  NR2 U24460 ( .I1(n18542), .I2(n18532), .O(n25195) );
  INV1S U24461 ( .I(n25195), .O(n25334) );
  NR2 U24462 ( .I1(n18543), .I2(n18533), .O(n25333) );
  MOAI1S U24463 ( .A1(n25334), .A2(n18829), .B1(n25333), .B2(n19719), .O(
        n18534) );
  ND2S U24464 ( .I1(n15891), .I2(n20534), .O(n18536) );
  ND2S U24465 ( .I1(n18536), .I2(n18535), .O(n15230) );
  INV1S U24466 ( .I(n29831), .O(n26445) );
  NR2 U24467 ( .I1(n18577), .I2(n18537), .O(n25217) );
  INV1S U24468 ( .I(n25217), .O(n25348) );
  NR2 U24469 ( .I1(n18579), .I2(n18538), .O(n25347) );
  MOAI1S U24470 ( .A1(n25348), .A2(n18829), .B1(n25347), .B2(n19719), .O(
        n18539) );
  ND2S U24471 ( .I1(n26445), .I2(n20562), .O(n18541) );
  ND2S U24472 ( .I1(n18541), .I2(n18540), .O(n15206) );
  NR2 U24473 ( .I1(n18542), .I2(n18577), .O(n25103) );
  INV1S U24474 ( .I(n25103), .O(n25358) );
  NR2 U24475 ( .I1(n18543), .I2(n18579), .O(n25356) );
  MOAI1S U24476 ( .A1(n25358), .A2(n18829), .B1(n25356), .B2(n19719), .O(
        n18544) );
  ND2S U24477 ( .I1(n26445), .I2(n20559), .O(n18546) );
  ND2S U24478 ( .I1(n18546), .I2(n18545), .O(n15214) );
  ND2S U24479 ( .I1(n15891), .I2(n20525), .O(n18548) );
  ND2S U24480 ( .I1(n18548), .I2(n18547), .O(n15126) );
  INV1S U24481 ( .I(n29831), .O(n26828) );
  INV1S U24482 ( .I(n25308), .O(n25342) );
  MOAI1S U24483 ( .A1(n25342), .A2(n18829), .B1(n25340), .B2(n19719), .O(
        n18549) );
  ND2S U24484 ( .I1(n26828), .I2(n20054), .O(n18551) );
  ND2S U24485 ( .I1(n18551), .I2(n18550), .O(n15222) );
  MUX2S U24486 ( .A(n30005), .B(n20156), .S(gray_img[1829]), .O(n18553) );
  ND2S U24487 ( .I1(n26828), .I2(n20156), .O(n18552) );
  ND2S U24488 ( .I1(n18553), .I2(n18552), .O(n15104) );
  ND2S U24489 ( .I1(n26445), .I2(n20368), .O(n18554) );
  ND2S U24490 ( .I1(n18555), .I2(n18554), .O(n15200) );
  ND2S U24491 ( .I1(n26445), .I2(n20379), .O(n18556) );
  ND2S U24492 ( .I1(n18557), .I2(n18556), .O(n15184) );
  ND2S U24493 ( .I1(n25389), .I2(n20054), .O(n18559) );
  ND2S U24494 ( .I1(n25389), .I2(n20063), .O(n18561) );
  MUX2S U24495 ( .A(n30005), .B(n20063), .S(gray_img[1910]), .O(n18560) );
  ND2S U24496 ( .I1(n18561), .I2(n18560), .O(n15290) );
  ND2S U24497 ( .I1(n25444), .I2(n20525), .O(n18563) );
  ND2S U24498 ( .I1(n25389), .I2(n20562), .O(n18565) );
  NR2 U24499 ( .I1(n18572), .I2(n18567), .O(n25286) );
  MOAI1S U24500 ( .A1(n20322), .A2(n25287), .B1(n25193), .B2(n25286), .O(
        n18568) );
  MUX2S U24501 ( .A(n15904), .B(n20843), .S(gray_img[1317]), .O(n18570) );
  ND2S U24502 ( .I1(n15891), .I2(n20843), .O(n18569) );
  ND2S U24503 ( .I1(n18570), .I2(n18569), .O(n15168) );
  NR2 U24504 ( .I1(n18572), .I2(n18578), .O(n25292) );
  MOAI1S U24505 ( .A1(n20322), .A2(n25293), .B1(n25193), .B2(n25292), .O(
        n18573) );
  ND2S U24506 ( .I1(n26445), .I2(n20811), .O(n18574) );
  ND2S U24507 ( .I1(n18575), .I2(n18574), .O(n15152) );
  NR2 U24508 ( .I1(n18577), .I2(n18576), .O(n19788) );
  NR2 U24509 ( .I1(n18579), .I2(n18578), .O(n25061) );
  AOI22S U24510 ( .A1(n19788), .A2(n19720), .B1(n25061), .B2(n19719), .O(
        n25943) );
  ND2S U24511 ( .I1(n15891), .I2(n25942), .O(n18581) );
  MUX2S U24512 ( .A(n30005), .B(n25942), .S(gray_img[2037]), .O(n18580) );
  ND2S U24513 ( .I1(n18581), .I2(n18580), .O(n15078) );
  MUX2S U24514 ( .A(n30005), .B(n25942), .S(gray_img[2035]), .O(n18582) );
  ND2S U24515 ( .I1(n18583), .I2(n18582), .O(n14679) );
  MUX2S U24516 ( .A(n30005), .B(n25942), .S(gray_img[2033]), .O(n18584) );
  ND2S U24517 ( .I1(n18585), .I2(n18584), .O(n14278) );
  MOAI1S U24518 ( .A1(n18829), .A2(n25297), .B1(n19719), .B2(n25296), .O(
        n18586) );
  ND2S U24519 ( .I1(n25389), .I2(n20725), .O(n18588) );
  INV1S U24520 ( .I(n27447), .O(n20808) );
  MOAI1S U24521 ( .A1(n18829), .A2(n25301), .B1(n19719), .B2(n25300), .O(
        n18589) );
  ND2S U24522 ( .I1(n25444), .I2(n20124), .O(n18591) );
  ND2S U24523 ( .I1(n26445), .I2(n20725), .O(n18593) );
  ND2S U24524 ( .I1(n18593), .I2(n18592), .O(n15174) );
  ND2S U24525 ( .I1(n15891), .I2(n20124), .O(n18595) );
  ND2S U24526 ( .I1(n18595), .I2(n18594), .O(n15190) );
  INV1S U24527 ( .I(n25086), .O(n18625) );
  MOAI1S U24528 ( .A1(n18625), .A2(n25287), .B1(n25085), .B2(n25286), .O(
        n18596) );
  MUX2S U24529 ( .A(n30005), .B(n20129), .S(gray_img[1309]), .O(n18598) );
  ND2S U24530 ( .I1(n27751), .I2(n20129), .O(n18597) );
  ND2S U24531 ( .I1(n18598), .I2(n18597), .O(n15169) );
  MOAI1S U24532 ( .A1(n18625), .A2(n25293), .B1(n25085), .B2(n25292), .O(
        n18599) );
  ND2S U24533 ( .I1(n27751), .I2(n20293), .O(n18600) );
  ND2S U24534 ( .I1(n18601), .I2(n18600), .O(n15153) );
  MOAI1S U24535 ( .A1(n18625), .A2(n25058), .B1(n25085), .B2(n25057), .O(
        n18602) );
  MUX2S U24536 ( .A(n30005), .B(n20599), .S(gray_img[1693]), .O(n18604) );
  ND2S U24537 ( .I1(n26445), .I2(n20599), .O(n18603) );
  ND2S U24538 ( .I1(n18604), .I2(n18603), .O(n15121) );
  MOAI1S U24539 ( .A1(n18625), .A2(n25054), .B1(n25085), .B2(n25053), .O(
        n18605) );
  MUX2S U24540 ( .A(n30005), .B(n20596), .S(gray_img[1565]), .O(n18607) );
  ND2S U24541 ( .I1(n26445), .I2(n20596), .O(n18606) );
  ND2S U24542 ( .I1(n18607), .I2(n18606), .O(n15137) );
  INV1S U24543 ( .I(n19788), .O(n25062) );
  MOAI1S U24544 ( .A1(n18625), .A2(n25062), .B1(n25085), .B2(n25061), .O(
        n18608) );
  ND2S U24545 ( .I1(n15890), .I2(n19970), .O(n18609) );
  ND2S U24546 ( .I1(n18610), .I2(n18609), .O(n15285) );
  MOAI1S U24547 ( .A1(n18625), .A2(n25297), .B1(n25085), .B2(n25296), .O(
        n18611) );
  ND2S U24548 ( .I1(n27751), .I2(n20159), .O(n18612) );
  ND2S U24549 ( .I1(n18613), .I2(n18612), .O(n15185) );
  ND2S U24550 ( .I1(n15890), .I2(n20596), .O(n18614) );
  ND2S U24551 ( .I1(n18615), .I2(n18614), .O(n15333) );
  MOAI1S U24552 ( .A1(n18625), .A2(n25301), .B1(n25085), .B2(n25300), .O(
        n18616) );
  ND2S U24553 ( .I1(n15891), .I2(n20184), .O(n18617) );
  ND2S U24554 ( .I1(n18618), .I2(n18617), .O(n15201) );
  INV1S U24555 ( .I(n29825), .O(n25389) );
  ND2S U24556 ( .I1(n25389), .I2(n20159), .O(n18619) );
  ND2S U24557 ( .I1(n18620), .I2(n18619), .O(n15381) );
  MUX2S U24558 ( .A(n30005), .B(n20129), .S(gray_img[1305]), .O(n18622) );
  ND2S U24559 ( .I1(n18622), .I2(n18621), .O(n14369) );
  ND2S U24560 ( .I1(n25389), .I2(n20184), .O(n18623) );
  ND2S U24561 ( .I1(n18624), .I2(n18623), .O(n15397) );
  MOAI1S U24562 ( .A1(n18625), .A2(n25066), .B1(n25085), .B2(n25065), .O(
        n18626) );
  ND2S U24563 ( .I1(n27751), .I2(n20296), .O(n18627) );
  ND2S U24564 ( .I1(n18628), .I2(n18627), .O(n15105) );
  ND2S U24565 ( .I1(n18630), .I2(n18629), .O(n14754) );
  ND2S U24566 ( .I1(n18632), .I2(n18631), .O(n14554) );
  ND2S U24567 ( .I1(n15891), .I2(n19970), .O(n18633) );
  ND2S U24568 ( .I1(n18634), .I2(n18633), .O(n15089) );
  ND2S U24569 ( .I1(n18636), .I2(n18635), .O(n14786) );
  ND2S U24570 ( .I1(n18638), .I2(n18637), .O(n14586) );
  ND2S U24571 ( .I1(n18640), .I2(n18639), .O(n14385) );
  INV1S U24572 ( .I(n25273), .O(n25254) );
  NR2 U24573 ( .I1(n18820), .I2(n24996), .O(n19407) );
  INV1S U24574 ( .I(n19407), .O(n18789) );
  MOAI1S U24575 ( .A1(n25254), .A2(n18789), .B1(n25271), .B2(n19406), .O(
        n18643) );
  ND2S U24576 ( .I1(n15891), .I2(n20082), .O(n18645) );
  ND2S U24577 ( .I1(n18645), .I2(n18644), .O(n15261) );
  ND2S U24578 ( .I1(n15890), .I2(n20082), .O(n18647) );
  ND2S U24579 ( .I1(n18647), .I2(n18646), .O(n15457) );
  MOAI1S U24580 ( .A1(n25342), .A2(n18789), .B1(n25340), .B2(n19406), .O(
        n18648) );
  ND2S U24581 ( .I1(n15891), .I2(n20568), .O(n18650) );
  INV1S U24582 ( .I(n27447), .O(n25928) );
  ND2S U24583 ( .I1(n18650), .I2(n18649), .O(n15221) );
  MOAI1S U24584 ( .A1(n25362), .A2(n18789), .B1(n25361), .B2(n19406), .O(
        n18651) );
  ND2S U24585 ( .I1(n27751), .I2(n20486), .O(n18653) );
  ND2S U24586 ( .I1(n18653), .I2(n18652), .O(n15245) );
  MOAI1S U24587 ( .A1(n25358), .A2(n18789), .B1(n25356), .B2(n19406), .O(
        n18654) );
  ND2S U24588 ( .I1(n26445), .I2(n20452), .O(n18656) );
  ND2S U24589 ( .I1(n18656), .I2(n18655), .O(n15213) );
  MOAI1S U24590 ( .A1(n25334), .A2(n18789), .B1(n25333), .B2(n19406), .O(
        n18657) );
  ND2S U24591 ( .I1(n15891), .I2(n20565), .O(n18659) );
  ND2S U24592 ( .I1(n18659), .I2(n18658), .O(n15229) );
  MOAI1S U24593 ( .A1(n25348), .A2(n18789), .B1(n25347), .B2(n19406), .O(
        n18660) );
  ND2S U24594 ( .I1(n26828), .I2(n20099), .O(n18662) );
  ND2S U24595 ( .I1(n18662), .I2(n18661), .O(n15205) );
  INV1S U24596 ( .I(n27447), .O(n20830) );
  NR2 U24597 ( .I1(n18883), .I2(n18820), .O(n25373) );
  INV1S U24598 ( .I(n25373), .O(n18689) );
  MOAI1S U24599 ( .A1(n18689), .A2(n25054), .B1(n25371), .B2(n25053), .O(
        n18663) );
  ND2S U24600 ( .I1(n27751), .I2(n20839), .O(n18664) );
  ND2S U24601 ( .I1(n18665), .I2(n18664), .O(n15134) );
  MOAI1S U24602 ( .A1(n18689), .A2(n25293), .B1(n25371), .B2(n25292), .O(
        n18666) );
  ND2S U24603 ( .I1(n26445), .I2(n20821), .O(n18667) );
  ND2S U24604 ( .I1(n18668), .I2(n18667), .O(n15150) );
  MOAI1S U24605 ( .A1(n18689), .A2(n25297), .B1(n25371), .B2(n25296), .O(
        n18669) );
  ND2S U24606 ( .I1(n26828), .I2(n20857), .O(n18670) );
  ND2S U24607 ( .I1(n18671), .I2(n18670), .O(n15182) );
  ND2S U24608 ( .I1(n25389), .I2(n20099), .O(n18673) );
  MOAI1S U24609 ( .A1(n18689), .A2(n25287), .B1(n25371), .B2(n25286), .O(
        n18674) );
  ND2S U24610 ( .I1(n15891), .I2(n20833), .O(n18675) );
  ND2S U24611 ( .I1(n18676), .I2(n18675), .O(n15166) );
  MOAI1S U24612 ( .A1(n18689), .A2(n25301), .B1(n25371), .B2(n25300), .O(
        n18677) );
  ND2S U24613 ( .I1(n26828), .I2(n20854), .O(n18678) );
  ND2S U24614 ( .I1(n18679), .I2(n18678), .O(n15198) );
  MOAI1S U24615 ( .A1(n18689), .A2(n25066), .B1(n25371), .B2(n25065), .O(
        n18680) );
  ND2S U24616 ( .I1(n15891), .I2(n20862), .O(n18681) );
  ND2S U24617 ( .I1(n18682), .I2(n18681), .O(n15102) );
  MOAI1S U24618 ( .A1(n18689), .A2(n25058), .B1(n25371), .B2(n25057), .O(
        n18683) );
  ND2S U24619 ( .I1(n26445), .I2(n20846), .O(n18684) );
  ND2S U24620 ( .I1(n18685), .I2(n18684), .O(n15118) );
  INV1S U24621 ( .I(n25246), .O(n25258) );
  MOAI1S U24622 ( .A1(n25258), .A2(n18789), .B1(n25257), .B2(n19406), .O(
        n18686) );
  ND2S U24623 ( .I1(n15891), .I2(n20496), .O(n18688) );
  ND2S U24624 ( .I1(n18688), .I2(n18687), .O(n15253) );
  MOAI1S U24625 ( .A1(n18689), .A2(n25062), .B1(n25371), .B2(n25061), .O(
        n18690) );
  ND2S U24626 ( .I1(n26445), .I2(n20849), .O(n18691) );
  ND2S U24627 ( .I1(n18692), .I2(n18691), .O(n15086) );
  MOAI1S U24628 ( .A1(n25367), .A2(n18789), .B1(n25370), .B2(n19406), .O(
        n18693) );
  ND2S U24629 ( .I1(n18695), .I2(n18694), .O(n14638) );
  ND2S U24630 ( .I1(n18697), .I2(n18696), .O(n14814) );
  ND2S U24631 ( .I1(n18699), .I2(n18698), .O(n14646) );
  ND2S U24632 ( .I1(n18701), .I2(n18700), .O(n14614) );
  NR2 U24633 ( .I1(n24997), .I2(n18819), .O(n25326) );
  INV1S U24634 ( .I(n25326), .O(n18812) );
  MOAI1S U24635 ( .A1(n18812), .A2(n25293), .B1(n25325), .B2(n25292), .O(
        n18702) );
  ND2S U24636 ( .I1(n27751), .I2(n20035), .O(n18704) );
  INV1S U24637 ( .I(n27447), .O(n20842) );
  ND2S U24638 ( .I1(n18704), .I2(n18703), .O(n15155) );
  MOAI1S U24639 ( .A1(n18812), .A2(n25287), .B1(n25325), .B2(n25286), .O(
        n18705) );
  ND2S U24640 ( .I1(n27751), .I2(n20427), .O(n18707) );
  ND2S U24641 ( .I1(n18707), .I2(n18706), .O(n15171) );
  MOAI1S U24642 ( .A1(n18812), .A2(n25054), .B1(n25325), .B2(n25053), .O(
        n18708) );
  ND2S U24643 ( .I1(n26828), .I2(n20550), .O(n18710) );
  ND2S U24644 ( .I1(n18710), .I2(n18709), .O(n15139) );
  ND2S U24645 ( .I1(n18712), .I2(n18711), .O(n14654) );
  MOAI1S U24646 ( .A1(n18812), .A2(n25058), .B1(n25325), .B2(n25057), .O(
        n18713) );
  ND2S U24647 ( .I1(n26828), .I2(n20531), .O(n18715) );
  ND2S U24648 ( .I1(n18715), .I2(n18714), .O(n15123) );
  ND2S U24649 ( .I1(n15890), .I2(n20550), .O(n18717) );
  ND2S U24650 ( .I1(n18717), .I2(n18716), .O(n15335) );
  MOAI1S U24651 ( .A1(n18812), .A2(n25297), .B1(n25325), .B2(n25296), .O(
        n18718) );
  ND2S U24652 ( .I1(n26828), .I2(n20553), .O(n18720) );
  ND2S U24653 ( .I1(n18720), .I2(n18719), .O(n15187) );
  ND2S U24654 ( .I1(n18722), .I2(n18721), .O(n14355) );
  ND2S U24655 ( .I1(n18724), .I2(n18723), .O(n14556) );
  ND2S U24656 ( .I1(n18726), .I2(n18725), .O(n14756) );
  ND2S U24657 ( .I1(n18728), .I2(n18727), .O(n14371) );
  MUX2S U24658 ( .A(n20842), .B(n20427), .S(gray_img[1290]), .O(n18729) );
  ND2S U24659 ( .I1(n18730), .I2(n18729), .O(n14572) );
  ND2S U24660 ( .I1(n18732), .I2(n18731), .O(n14772) );
  INV1S U24661 ( .I(medfilt_out_reg[0]), .O(n18735) );
  OAI12HS U24662 ( .B1(n18735), .B2(n18734), .A1(n18733), .O(n19092) );
  MOAI1S U24663 ( .A1(n18789), .A2(n25293), .B1(n19406), .B2(n25292), .O(
        n18736) );
  ND2S U24664 ( .I1(n19092), .I2(n20556), .O(n18738) );
  ND2S U24665 ( .I1(n18738), .I2(n18737), .O(n13928) );
  INV1S U24666 ( .I(n25245), .O(n18774) );
  MOAI1S U24667 ( .A1(n18774), .A2(n25066), .B1(n25244), .B2(n25065), .O(
        n18739) );
  MUX2S U24668 ( .A(n30005), .B(n20142), .S(gray_img[1837]), .O(n18741) );
  ND2S U24669 ( .I1(n26828), .I2(n20142), .O(n18740) );
  ND2S U24670 ( .I1(n18741), .I2(n18740), .O(n15103) );
  MOAI1S U24671 ( .A1(n18789), .A2(n25066), .B1(n19406), .B2(n25065), .O(
        n18742) );
  ND2S U24672 ( .I1(n19092), .I2(n20430), .O(n18744) );
  ND2S U24673 ( .I1(n18744), .I2(n18743), .O(n13844) );
  ND2S U24674 ( .I1(n15891), .I2(n20556), .O(n18746) );
  ND2S U24675 ( .I1(n18746), .I2(n18745), .O(n15141) );
  MOAI1S U24676 ( .A1(n18789), .A2(n25287), .B1(n19406), .B2(n25286), .O(
        n18747) );
  ND2S U24677 ( .I1(n15891), .I2(n20571), .O(n18749) );
  ND2S U24678 ( .I1(n18749), .I2(n18748), .O(n15157) );
  ND2S U24679 ( .I1(n15891), .I2(n20430), .O(n18751) );
  ND2S U24680 ( .I1(n18751), .I2(n18750), .O(n15093) );
  MOAI1S U24681 ( .A1(n18774), .A2(n25062), .B1(n25244), .B2(n25061), .O(
        n18752) );
  MUX2S U24682 ( .A(n30005), .B(n20202), .S(gray_img[1965]), .O(n18754) );
  ND2S U24683 ( .I1(n26828), .I2(n20202), .O(n18753) );
  ND2S U24684 ( .I1(n18754), .I2(n18753), .O(n15087) );
  ND2S U24685 ( .I1(n25444), .I2(n20571), .O(n18756) );
  ND2S U24686 ( .I1(n18756), .I2(n18755), .O(n15353) );
  MOAI1S U24687 ( .A1(n18774), .A2(n25058), .B1(n25244), .B2(n25057), .O(
        n18757) );
  ND2S U24688 ( .I1(n15891), .I2(n20827), .O(n18758) );
  ND2S U24689 ( .I1(n18759), .I2(n18758), .O(n15119) );
  MOAI1S U24690 ( .A1(n18774), .A2(n25054), .B1(n25244), .B2(n25053), .O(
        n18760) );
  ND2S U24691 ( .I1(n27751), .I2(n20395), .O(n18761) );
  ND2S U24692 ( .I1(n18762), .I2(n18761), .O(n15135) );
  MOAI1S U24693 ( .A1(n18789), .A2(n25054), .B1(n19406), .B2(n25053), .O(
        n18763) );
  ND2S U24694 ( .I1(n27751), .I2(n20509), .O(n18765) );
  ND2S U24695 ( .I1(n18765), .I2(n18764), .O(n15125) );
  MUX2S U24696 ( .A(n30005), .B(n20142), .S(gray_img[1835]), .O(n18767) );
  ND2S U24697 ( .I1(n18767), .I2(n18766), .O(n14704) );
  MOAI1S U24698 ( .A1(n18789), .A2(n25297), .B1(n19406), .B2(n25296), .O(
        n18768) );
  ND2S U24699 ( .I1(n19092), .I2(n20655), .O(n18770) );
  ND2S U24700 ( .I1(n18770), .I2(n18769), .O(n14010) );
  MOAI1S U24701 ( .A1(n18774), .A2(n25293), .B1(n25244), .B2(n25292), .O(
        n18771) );
  MUX2S U24702 ( .A(n30005), .B(n20814), .S(gray_img[1453]), .O(n18773) );
  ND2S U24703 ( .I1(n15891), .I2(n20814), .O(n18772) );
  ND2S U24704 ( .I1(n18773), .I2(n18772), .O(n15151) );
  MOAI1S U24705 ( .A1(n18774), .A2(n25287), .B1(n25244), .B2(n25286), .O(
        n18775) );
  ND2S U24706 ( .I1(n27751), .I2(n20836), .O(n18776) );
  ND2S U24707 ( .I1(n18777), .I2(n18776), .O(n15167) );
  MOAI1S U24708 ( .A1(n18789), .A2(n25301), .B1(n19406), .B2(n25300), .O(
        n18778) );
  ND2S U24709 ( .I1(n19092), .I2(n20716), .O(n18780) );
  ND2S U24710 ( .I1(n18780), .I2(n18779), .O(n14075) );
  ND2S U24711 ( .I1(n18782), .I2(n18781), .O(n14504) );
  MUX2S U24712 ( .A(n30005), .B(n20202), .S(gray_img[1961]), .O(n18784) );
  ND2S U24713 ( .I1(n18784), .I2(n18783), .O(n14287) );
  ND2S U24714 ( .I1(n18786), .I2(n18785), .O(n14293) );
  ND2S U24715 ( .I1(n18788), .I2(n18787), .O(n14694) );
  MOAI1S U24716 ( .A1(n18789), .A2(n25058), .B1(n19406), .B2(n25057), .O(
        n18790) );
  MUX2S U24717 ( .A(n29032), .B(n20547), .S(gray_img[1785]), .O(n18791) );
  ND2S U24718 ( .I1(n18792), .I2(n18791), .O(n14309) );
  ND2S U24719 ( .I1(n18794), .I2(n18793), .O(n14710) );
  ND2S U24720 ( .I1(n18796), .I2(n18795), .O(n14325) );
  ND2S U24721 ( .I1(n18798), .I2(n18797), .O(n14726) );
  ND2S U24722 ( .I1(n26445), .I2(n20655), .O(n18800) );
  ND2S U24723 ( .I1(n18800), .I2(n18799), .O(n15173) );
  ND2S U24724 ( .I1(n18802), .I2(n18801), .O(n14289) );
  ND2S U24725 ( .I1(n15891), .I2(n20716), .O(n18804) );
  ND2S U24726 ( .I1(n18804), .I2(n18803), .O(n15189) );
  ND2S U24727 ( .I1(n15891), .I2(n20547), .O(n18806) );
  ND2S U24728 ( .I1(n18806), .I2(n18805), .O(n15109) );
  ND2S U24729 ( .I1(n27751), .I2(n20472), .O(n18808) );
  ND2S U24730 ( .I1(n18808), .I2(n18807), .O(n15237) );
  MOAI1S U24731 ( .A1(n18812), .A2(n25062), .B1(n25325), .B2(n25061), .O(
        n18809) );
  ND2S U24732 ( .I1(n26445), .I2(n20424), .O(n18811) );
  ND2S U24733 ( .I1(n18811), .I2(n18810), .O(n15091) );
  MOAI1S U24734 ( .A1(n18812), .A2(n25066), .B1(n25325), .B2(n25065), .O(
        n18813) );
  ND2S U24735 ( .I1(n27751), .I2(n20319), .O(n18815) );
  ND2S U24736 ( .I1(n18815), .I2(n18814), .O(n15107) );
  MOAI1S U24737 ( .A1(n18829), .A2(n25293), .B1(n19719), .B2(n25292), .O(
        n18816) );
  ND2S U24738 ( .I1(n26445), .I2(n20512), .O(n18818) );
  ND2S U24739 ( .I1(n18818), .I2(n18817), .O(n15142) );
  NR2 U24740 ( .I1(n18820), .I2(n18819), .O(n25283) );
  INV1S U24741 ( .I(n25283), .O(n18854) );
  MOAI1S U24742 ( .A1(n18854), .A2(n25287), .B1(n25282), .B2(n25286), .O(
        n18823) );
  ND2S U24743 ( .I1(n15891), .I2(n20695), .O(n18825) );
  ND2S U24744 ( .I1(n18825), .I2(n18824), .O(n15165) );
  MOAI1S U24745 ( .A1(n18854), .A2(n25293), .B1(n25282), .B2(n25292), .O(
        n18826) );
  ND2S U24746 ( .I1(n15891), .I2(n20709), .O(n18828) );
  ND2S U24747 ( .I1(n18828), .I2(n18827), .O(n15149) );
  MOAI1S U24748 ( .A1(n18829), .A2(n25287), .B1(n19719), .B2(n25286), .O(
        n18830) );
  ND2S U24749 ( .I1(n15891), .I2(n20517), .O(n18832) );
  ND2S U24750 ( .I1(n18832), .I2(n18831), .O(n15158) );
  MOAI1S U24751 ( .A1(n18854), .A2(n25058), .B1(n25282), .B2(n25057), .O(
        n18833) );
  ND2S U24752 ( .I1(n27751), .I2(n20737), .O(n18835) );
  ND2S U24753 ( .I1(n18835), .I2(n18834), .O(n15117) );
  MOAI1S U24754 ( .A1(n18854), .A2(n25054), .B1(n25282), .B2(n25053), .O(
        n18836) );
  ND2S U24755 ( .I1(n26828), .I2(n20731), .O(n18838) );
  ND2S U24756 ( .I1(n18838), .I2(n18837), .O(n15133) );
  ND2S U24757 ( .I1(n18840), .I2(n18839), .O(n14291) );
  ND2S U24758 ( .I1(n18842), .I2(n18841), .O(n14662) );
  ND2S U24759 ( .I1(n18844), .I2(n18843), .O(n14307) );
  INV1S U24760 ( .I(n25218), .O(n20865) );
  MOAI1S U24761 ( .A1(n20865), .A2(n25058), .B1(n25216), .B2(n25057), .O(
        n18845) );
  ND2S U24762 ( .I1(n26445), .I2(n20583), .O(n18846) );
  ND2S U24763 ( .I1(n18847), .I2(n18846), .O(n15124) );
  MOAI1S U24764 ( .A1(n20865), .A2(n25066), .B1(n25216), .B2(n25065), .O(
        n18848) );
  MUX2S U24765 ( .A(n29032), .B(n20376), .S(gray_img[1797]), .O(n18850) );
  ND2S U24766 ( .I1(n26828), .I2(n20376), .O(n18849) );
  ND2S U24767 ( .I1(n18850), .I2(n18849), .O(n15108) );
  MOAI1S U24768 ( .A1(n18854), .A2(n25066), .B1(n25282), .B2(n25065), .O(
        n18851) );
  ND2S U24769 ( .I1(n15891), .I2(n20740), .O(n18853) );
  ND2S U24770 ( .I1(n18853), .I2(n18852), .O(n15101) );
  MOAI1S U24771 ( .A1(n18854), .A2(n25062), .B1(n25282), .B2(n25061), .O(
        n18855) );
  ND2S U24772 ( .I1(n26828), .I2(n20746), .O(n18857) );
  ND2S U24773 ( .I1(n18857), .I2(n18856), .O(n15085) );
  MOAI1S U24774 ( .A1(n20865), .A2(n25293), .B1(n25216), .B2(n25292), .O(
        n18858) );
  MUX2S U24775 ( .A(n30005), .B(n20359), .S(gray_img[1413]), .O(n18860) );
  ND2S U24776 ( .I1(n15891), .I2(n20359), .O(n18859) );
  ND2S U24777 ( .I1(n18860), .I2(n18859), .O(n15156) );
  MOAI1S U24778 ( .A1(n20865), .A2(n25287), .B1(n25216), .B2(n25286), .O(
        n18861) );
  ND2S U24779 ( .I1(n26828), .I2(n20392), .O(n18862) );
  ND2S U24780 ( .I1(n18863), .I2(n18862), .O(n15172) );
  ND2S U24781 ( .I1(n18865), .I2(n18864), .O(n14557) );
  MUX2S U24782 ( .A(n30005), .B(n20359), .S(gray_img[1409]), .O(n18867) );
  ND2S U24783 ( .I1(n18867), .I2(n18866), .O(n14356) );
  MUX2S U24784 ( .A(n30005), .B(n20359), .S(gray_img[1411]), .O(n18869) );
  ND2S U24785 ( .I1(n18869), .I2(n18868), .O(n14757) );
  ND2S U24786 ( .I1(n18871), .I2(n18870), .O(n14573) );
  ND2S U24787 ( .I1(n18873), .I2(n18872), .O(n14773) );
  ND2S U24788 ( .I1(n18875), .I2(n18874), .O(n14372) );
  ND2S U24789 ( .I1(n18877), .I2(n18876), .O(n14308) );
  MOAI1S U24790 ( .A1(n20865), .A2(n25062), .B1(n25216), .B2(n25061), .O(
        n18878) );
  ND2S U24791 ( .I1(n15891), .I2(n20373), .O(n18879) );
  ND2S U24792 ( .I1(n18880), .I2(n18879), .O(n15092) );
  ND2S U24793 ( .I1(n18882), .I2(n18881), .O(n14292) );
  NR2 U24794 ( .I1(n18883), .I2(n24972), .O(n25274) );
  INV1S U24795 ( .I(n25274), .O(n20334) );
  MOAI1S U24796 ( .A1(n20334), .A2(n25293), .B1(n25272), .B2(n25292), .O(
        n18885) );
  ND2S U24797 ( .I1(n27751), .I2(n20193), .O(n18886) );
  ND2S U24798 ( .I1(n18887), .I2(n18886), .O(n15154) );
  MOAI1S U24799 ( .A1(n20334), .A2(n25287), .B1(n25272), .B2(n25286), .O(
        n18888) );
  ND2S U24800 ( .I1(n27751), .I2(n20362), .O(n18889) );
  ND2S U24801 ( .I1(n18890), .I2(n18889), .O(n15170) );
  ND2S U24802 ( .I1(n15890), .I2(n20193), .O(n18891) );
  MOAI1S U24803 ( .A1(n20334), .A2(n25058), .B1(n25272), .B2(n25057), .O(
        n18893) );
  ND2S U24804 ( .I1(n26445), .I2(n20605), .O(n18894) );
  ND2S U24805 ( .I1(n18895), .I2(n18894), .O(n15122) );
  MOAI1S U24806 ( .A1(n20334), .A2(n25054), .B1(n25272), .B2(n25053), .O(
        n18896) );
  ND2S U24807 ( .I1(n26445), .I2(n20602), .O(n18897) );
  ND2S U24808 ( .I1(n18898), .I2(n18897), .O(n15138) );
  MOAI1S U24809 ( .A1(n20334), .A2(n25062), .B1(n25272), .B2(n25061), .O(
        n18899) );
  ND2S U24810 ( .I1(n15891), .I2(n20389), .O(n18900) );
  ND2S U24811 ( .I1(n18901), .I2(n18900), .O(n15090) );
  ND2S U24812 ( .I1(n18903), .I2(n18902), .O(n14290) );
  NR2 U24813 ( .I1(n25050), .I2(n24996), .O(n19845) );
  INV1S U24814 ( .I(n19845), .O(n18973) );
  MOAI1S U24815 ( .A1(n25358), .A2(n18973), .B1(n25356), .B2(n19844), .O(
        n18904) );
  MUX2S U24816 ( .A(n30005), .B(n20212), .S(gray_img[877]), .O(n18906) );
  ND2S U24817 ( .I1(n27751), .I2(n20212), .O(n18905) );
  ND2S U24818 ( .I1(n18906), .I2(n18905), .O(n15215) );
  MOAI1S U24819 ( .A1(n25342), .A2(n18973), .B1(n25340), .B2(n19844), .O(
        n18907) );
  MUX2S U24820 ( .A(n30005), .B(n20365), .S(gray_img[749]), .O(n18909) );
  ND2S U24821 ( .I1(n26828), .I2(n20365), .O(n18908) );
  ND2S U24822 ( .I1(n18909), .I2(n18908), .O(n15223) );
  MOAI1S U24823 ( .A1(n25348), .A2(n18973), .B1(n25347), .B2(n19844), .O(
        n18910) );
  MUX2S U24824 ( .A(n30005), .B(n20384), .S(gray_img[1005]), .O(n18912) );
  ND2S U24825 ( .I1(n26445), .I2(n20384), .O(n18911) );
  ND2S U24826 ( .I1(n18912), .I2(n18911), .O(n15207) );
  ND2S U24827 ( .I1(n25389), .I2(n20212), .O(n18913) );
  ND2S U24828 ( .I1(n18916), .I2(n18915), .O(n14415) );
  ND2S U24829 ( .I1(n18918), .I2(n18917), .O(n14423) );
  ND2S U24830 ( .I1(n18920), .I2(n18919), .O(n14624) );
  MUX2S U24831 ( .A(n25928), .B(n20384), .S(gray_img[1001]), .O(n18922) );
  ND2S U24832 ( .I1(n18922), .I2(n18921), .O(n14407) );
  NR2 U24833 ( .I1(n24997), .I2(n25049), .O(n19914) );
  INV1S U24834 ( .I(n19914), .O(n19001) );
  MOAI1S U24835 ( .A1(n25334), .A2(n19001), .B1(n25333), .B2(n19913), .O(
        n18923) );
  ND2S U24836 ( .I1(n26445), .I2(n20591), .O(n18924) );
  ND2S U24837 ( .I1(n18925), .I2(n18924), .O(n15236) );
  MOAI1S U24838 ( .A1(n25362), .A2(n19001), .B1(n25361), .B2(n19913), .O(
        n18926) );
  MUX2S U24839 ( .A(n30005), .B(n20147), .S(gray_img[325]), .O(n18928) );
  ND2S U24840 ( .I1(n15891), .I2(n20147), .O(n18927) );
  ND2S U24841 ( .I1(n18928), .I2(n18927), .O(n15252) );
  MOAI1S U24842 ( .A1(n25348), .A2(n19001), .B1(n25347), .B2(n19913), .O(
        n18929) );
  ND2S U24843 ( .I1(n26445), .I2(n20580), .O(n18930) );
  ND2S U24844 ( .I1(n18931), .I2(n18930), .O(n15212) );
  ND2S U24845 ( .I1(n25389), .I2(n20580), .O(n18932) );
  ND2S U24846 ( .I1(n18933), .I2(n18932), .O(n15408) );
  ND2S U24847 ( .I1(n25389), .I2(n20147), .O(n18934) );
  MOAI1S U24848 ( .A1(n25062), .A2(n19001), .B1(n25061), .B2(n19913), .O(
        n18936) );
  MUX2S U24849 ( .A(n30056), .B(n20209), .S(gray_img[1989]), .O(n18938) );
  ND2S U24850 ( .I1(n15891), .I2(n20209), .O(n18937) );
  ND2S U24851 ( .I1(n18938), .I2(n18937), .O(n15084) );
  ND2S U24852 ( .I1(n25389), .I2(n20209), .O(n18939) );
  ND2S U24853 ( .I1(n18942), .I2(n18941), .O(n14837) );
  ND2S U24854 ( .I1(n18944), .I2(n18943), .O(n14813) );
  MUX2S U24855 ( .A(n30056), .B(n20209), .S(gray_img[1986]), .O(n18946) );
  ND2S U24856 ( .I1(n18946), .I2(n18945), .O(n14485) );
  MUX2S U24857 ( .A(n29597), .B(n20209), .S(gray_img[1985]), .O(n18948) );
  ND2S U24858 ( .I1(n18948), .I2(n18947), .O(n14284) );
  MUX2S U24859 ( .A(n29566), .B(n20209), .S(gray_img[1987]), .O(n18950) );
  ND2S U24860 ( .I1(n18950), .I2(n18949), .O(n14685) );
  MOAI1S U24861 ( .A1(n18973), .A2(n25066), .B1(n19844), .B2(n25065), .O(
        n18951) );
  ND2S U24862 ( .I1(n15891), .I2(n20544), .O(n18953) );
  ND2S U24863 ( .I1(n18953), .I2(n18952), .O(n15095) );
  MOAI1S U24864 ( .A1(n18973), .A2(n25058), .B1(n19844), .B2(n25057), .O(
        n18954) );
  ND2S U24865 ( .I1(n26445), .I2(n20449), .O(n18956) );
  ND2S U24866 ( .I1(n18956), .I2(n18955), .O(n15111) );
  MOAI1S U24867 ( .A1(n18973), .A2(n25301), .B1(n19844), .B2(n25300), .O(
        n18957) );
  ND2S U24868 ( .I1(n26828), .I2(n20728), .O(n18959) );
  ND2S U24869 ( .I1(n18959), .I2(n18958), .O(n15191) );
  MOAI1S U24870 ( .A1(n18973), .A2(n25054), .B1(n19844), .B2(n25053), .O(
        n18960) );
  ND2S U24871 ( .I1(n27751), .I2(n20463), .O(n18962) );
  MUX2S U24872 ( .A(n30005), .B(n20463), .S(gray_img[1645]), .O(n18961) );
  ND2S U24873 ( .I1(n18962), .I2(n18961), .O(n15127) );
  ND2S U24874 ( .I1(n25389), .I2(n20728), .O(n18964) );
  ND2S U24875 ( .I1(n18964), .I2(n18963), .O(n15387) );
  MOAI1S U24876 ( .A1(n18973), .A2(n25297), .B1(n19844), .B2(n25296), .O(
        n18965) );
  ND2S U24877 ( .I1(n25444), .I2(n20719), .O(n18967) );
  ND2S U24878 ( .I1(n18967), .I2(n18966), .O(n15371) );
  MOAI1S U24879 ( .A1(n18973), .A2(n25287), .B1(n19844), .B2(n25286), .O(
        n18968) );
  ND2S U24880 ( .I1(n15891), .I2(n20722), .O(n18970) );
  ND2S U24881 ( .I1(n18970), .I2(n18969), .O(n15159) );
  ND2S U24882 ( .I1(n26445), .I2(n20719), .O(n18972) );
  ND2S U24883 ( .I1(n18972), .I2(n18971), .O(n15175) );
  MOAI1S U24884 ( .A1(n18973), .A2(n25293), .B1(n19844), .B2(n25292), .O(
        n18974) );
  ND2S U24885 ( .I1(n15891), .I2(n20440), .O(n18976) );
  ND2S U24886 ( .I1(n18976), .I2(n18975), .O(n15143) );
  MOAI1S U24887 ( .A1(n19001), .A2(n25066), .B1(n19913), .B2(n25065), .O(
        n18977) );
  ND2S U24888 ( .I1(n19092), .I2(n20504), .O(n18978) );
  ND2S U24889 ( .I1(n18979), .I2(n18978), .O(n13851) );
  MOAI1S U24890 ( .A1(n19001), .A2(n25054), .B1(n19913), .B2(n25053), .O(
        n18980) );
  ND2S U24891 ( .I1(n26828), .I2(n20528), .O(n18982) );
  ND2S U24892 ( .I1(n18982), .I2(n18981), .O(n15132) );
  ND2S U24893 ( .I1(n15891), .I2(n20504), .O(n18984) );
  ND2S U24894 ( .I1(n18984), .I2(n18983), .O(n15100) );
  MOAI1S U24895 ( .A1(n19001), .A2(n25058), .B1(n19913), .B2(n25057), .O(
        n18985) );
  ND2S U24896 ( .I1(n26828), .I2(n19955), .O(n18987) );
  ND2S U24897 ( .I1(n18987), .I2(n18986), .O(n15116) );
  MOAI1S U24898 ( .A1(n19001), .A2(n25287), .B1(n19913), .B2(n25286), .O(
        n18988) );
  ND2S U24899 ( .I1(n25389), .I2(n20734), .O(n18990) );
  ND2S U24900 ( .I1(n25389), .I2(n19955), .O(n18992) );
  ND2S U24901 ( .I1(n18992), .I2(n18991), .O(n15312) );
  ND2S U24902 ( .I1(n15890), .I2(n20528), .O(n18994) );
  ND2S U24903 ( .I1(n18994), .I2(n18993), .O(n15328) );
  MOAI1S U24904 ( .A1(n19001), .A2(n25301), .B1(n19913), .B2(n25300), .O(
        n18995) );
  ND2S U24905 ( .I1(n27751), .I2(n20743), .O(n18997) );
  ND2S U24906 ( .I1(n18997), .I2(n18996), .O(n15196) );
  MOAI1S U24907 ( .A1(n19001), .A2(n25293), .B1(n19913), .B2(n25292), .O(
        n18998) );
  ND2S U24908 ( .I1(n26828), .I2(n20684), .O(n19000) );
  ND2S U24909 ( .I1(n19000), .I2(n18999), .O(n15148) );
  MOAI1S U24910 ( .A1(n19001), .A2(n25297), .B1(n19913), .B2(n25296), .O(
        n19002) );
  ND2S U24911 ( .I1(n15891), .I2(n20702), .O(n19004) );
  ND2S U24912 ( .I1(n19004), .I2(n19003), .O(n15180) );
  ND2S U24913 ( .I1(n26828), .I2(n20734), .O(n19006) );
  ND2S U24914 ( .I1(n19006), .I2(n19005), .O(n15164) );
  MUX2S U24915 ( .A(n30005), .B(n20156), .S(gray_img[1824]), .O(n19008) );
  ND2S U24916 ( .I1(n15888), .I2(n20156), .O(n19007) );
  ND2S U24917 ( .I1(n19008), .I2(n19007), .O(n13855) );
  ND2S U24918 ( .I1(n15888), .I2(n20525), .O(n19009) );
  ND2S U24919 ( .I1(n19010), .I2(n19009), .O(n13909) );
  ND2S U24920 ( .I1(n15888), .I2(n20512), .O(n19011) );
  ND2S U24921 ( .I1(n19012), .I2(n19011), .O(n13929) );
  ND2S U24922 ( .I1(n15888), .I2(n20082), .O(n19013) );
  ND2S U24923 ( .I1(n19014), .I2(n19013), .O(n14259) );
  ND2S U24924 ( .I1(n15888), .I2(n20522), .O(n19015) );
  ND2S U24925 ( .I1(n19016), .I2(n19015), .O(n14216) );
  ND2S U24926 ( .I1(n15888), .I2(n20486), .O(n19017) );
  ND2S U24927 ( .I1(n19018), .I2(n19017), .O(n14215) );
  ND2S U24928 ( .I1(n15888), .I2(n20583), .O(n19019) );
  ND2S U24929 ( .I1(n19020), .I2(n19019), .O(n13907) );
  ND2S U24930 ( .I1(n15888), .I2(n20541), .O(n19021) );
  ND2S U24931 ( .I1(n19022), .I2(n19021), .O(n13865) );
  MUX2S U24932 ( .A(n30005), .B(n20147), .S(gray_img[320]), .O(n19024) );
  ND2S U24933 ( .I1(n15888), .I2(n20147), .O(n19023) );
  ND2S U24934 ( .I1(n19024), .I2(n19023), .O(n14222) );
  ND2S U24935 ( .I1(n15888), .I2(n19955), .O(n19025) );
  ND2S U24936 ( .I1(n19026), .I2(n19025), .O(n13883) );
  ND2S U24937 ( .I1(n15888), .I2(n20544), .O(n19027) );
  ND2S U24938 ( .I1(n19028), .I2(n19027), .O(n13846) );
  MUX2S U24939 ( .A(n30005), .B(n20202), .S(gray_img[1960]), .O(n19030) );
  ND2S U24940 ( .I1(n15888), .I2(n20202), .O(n19029) );
  ND2S U24941 ( .I1(n19030), .I2(n19029), .O(n13831) );
  ND2S U24942 ( .I1(n15888), .I2(n20580), .O(n19031) );
  ND2S U24943 ( .I1(n19032), .I2(n19031), .O(n14126) );
  ND2S U24944 ( .I1(n15888), .I2(n20599), .O(n19033) );
  ND2S U24945 ( .I1(n19034), .I2(n19033), .O(n13900) );
  ND2S U24946 ( .I1(n15888), .I2(n20821), .O(n19035) );
  ND2S U24947 ( .I1(n19036), .I2(n19035), .O(n13959) );
  ND2S U24948 ( .I1(n15888), .I2(n20496), .O(n19037) );
  ND2S U24949 ( .I1(n19038), .I2(n19037), .O(n14230) );
  ND2S U24950 ( .I1(n15888), .I2(n20142), .O(n19039) );
  ND2S U24951 ( .I1(n19040), .I2(n19039), .O(n13854) );
  ND2S U24952 ( .I1(n15888), .I2(n20734), .O(n19041) );
  ND2S U24953 ( .I1(n19042), .I2(n19041), .O(n13994) );
  MUX2S U24954 ( .A(n25928), .B(n20384), .S(gray_img[1000]), .O(n19044) );
  ND2S U24955 ( .I1(n15888), .I2(n20384), .O(n19043) );
  ND2S U24956 ( .I1(n19044), .I2(n19043), .O(n14107) );
  ND2S U24957 ( .I1(n15888), .I2(n20553), .O(n19045) );
  ND2S U24958 ( .I1(n19046), .I2(n19045), .O(n14073) );
  ND2S U24959 ( .I1(n15888), .I2(n20719), .O(n19047) );
  ND2S U24960 ( .I1(n19048), .I2(n19047), .O(n14019) );
  ND2S U24961 ( .I1(n15888), .I2(n20477), .O(n19049) );
  ND2S U24962 ( .I1(n19050), .I2(n19049), .O(n14187) );
  ND2S U24963 ( .I1(n15888), .I2(n20568), .O(n19051) );
  ND2S U24964 ( .I1(n19052), .I2(n19051), .O(n14142) );
  ND2S U24965 ( .I1(n15888), .I2(n20702), .O(n19053) );
  ND2S U24966 ( .I1(n19054), .I2(n19053), .O(n14038) );
  ND2S U24967 ( .I1(n15888), .I2(n20472), .O(n19055) );
  ND2S U24968 ( .I1(n19056), .I2(n19055), .O(n14186) );
  ND2S U24969 ( .I1(n15888), .I2(n20379), .O(n19057) );
  ND2S U24970 ( .I1(n19058), .I2(n19057), .O(n14056) );
  ND2S U24971 ( .I1(n15888), .I2(n20722), .O(n19059) );
  ND2S U24972 ( .I1(n19060), .I2(n19059), .O(n13989) );
  ND2S U24973 ( .I1(n15888), .I2(n20124), .O(n19061) );
  ND2S U24974 ( .I1(n19062), .I2(n19061), .O(n14076) );
  ND2S U24975 ( .I1(n15888), .I2(n20368), .O(n19063) );
  ND2S U24976 ( .I1(n19064), .I2(n19063), .O(n14086) );
  ND2S U24977 ( .I1(n15888), .I2(n20728), .O(n19065) );
  ND2S U24978 ( .I1(n19066), .I2(n19065), .O(n14077) );
  ND2S U24979 ( .I1(n15888), .I2(n20063), .O(n19067) );
  ND2S U24980 ( .I1(n19068), .I2(n19067), .O(n13845) );
  MUX2S U24981 ( .A(n30005), .B(n20565), .S(gray_img[632]), .O(n19070) );
  ND2S U24982 ( .I1(n15888), .I2(n20565), .O(n19069) );
  ND2S U24983 ( .I1(n19070), .I2(n19069), .O(n14171) );
  ND2S U24984 ( .I1(n15888), .I2(n20534), .O(n19071) );
  ND2S U24985 ( .I1(n19072), .I2(n19071), .O(n14172) );
  ND2S U24986 ( .I1(n15888), .I2(n20833), .O(n19073) );
  ND2S U24987 ( .I1(n19074), .I2(n19073), .O(n13996) );
  MUX2S U24988 ( .A(n30005), .B(n20452), .S(gray_img[888]), .O(n19076) );
  ND2S U24989 ( .I1(n15888), .I2(n20452), .O(n19075) );
  ND2S U24990 ( .I1(n19076), .I2(n19075), .O(n14127) );
  ND2S U24991 ( .I1(n15888), .I2(n20212), .O(n19077) );
  ND2S U24992 ( .I1(n19078), .I2(n19077), .O(n14129) );
  ND2S U24993 ( .I1(n15888), .I2(n20695), .O(n19079) );
  ND2S U24994 ( .I1(n19080), .I2(n19079), .O(n13995) );
  MUX2S U24995 ( .A(n30005), .B(n20099), .S(gray_img[1016]), .O(n19082) );
  ND2S U24996 ( .I1(n15888), .I2(n20099), .O(n19081) );
  ND2S U24997 ( .I1(n19082), .I2(n19081), .O(n14098) );
  ND2S U24998 ( .I1(n15888), .I2(n20547), .O(n19084) );
  ND2S U24999 ( .I1(n19084), .I2(n19083), .O(n13864) );
  ND2S U25000 ( .I1(n15888), .I2(n20571), .O(n19086) );
  ND2S U25001 ( .I1(n19086), .I2(n19085), .O(n13987) );
  INV1S U25002 ( .I(n24925), .O(n24930) );
  AOI22S U25003 ( .A1(n24069), .A2(n19089), .B1(n24930), .B2(n19088), .O(
        n19090) );
  ND2S U25004 ( .I1(n19091), .I2(n19090), .O(n15807) );
  ND2S U25005 ( .I1(n15888), .I2(n20293), .O(n19093) );
  ND2S U25006 ( .I1(n19094), .I2(n19093), .O(n13976) );
  MUX2S U25007 ( .A(n29032), .B(n20184), .S(gray_img[1048]), .O(n19096) );
  ND2S U25008 ( .I1(n15888), .I2(n20184), .O(n19095) );
  ND2S U25009 ( .I1(n19096), .I2(n19095), .O(n14087) );
  ND2S U25010 ( .I1(n15888), .I2(n20854), .O(n19097) );
  ND2S U25011 ( .I1(n19098), .I2(n19097), .O(n14084) );
  ND2S U25012 ( .I1(n15888), .I2(n20159), .O(n19099) );
  ND2S U25013 ( .I1(n19100), .I2(n19099), .O(n14064) );
  ND2S U25014 ( .I1(n15888), .I2(n20839), .O(n19101) );
  ND2S U25015 ( .I1(n19102), .I2(n19101), .O(n13917) );
  ND2S U25016 ( .I1(n15888), .I2(n20737), .O(n19103) );
  ND2S U25017 ( .I1(n19104), .I2(n19103), .O(n13888) );
  ND2S U25018 ( .I1(n15888), .I2(n20373), .O(n19105) );
  ND2S U25019 ( .I1(n19106), .I2(n19105), .O(n13843) );
  ND2S U25020 ( .I1(n15888), .I2(n20362), .O(n19107) );
  ND2S U25021 ( .I1(n19108), .I2(n19107), .O(n14000) );
  MUX2S U25022 ( .A(n30005), .B(n20359), .S(gray_img[1408]), .O(n19110) );
  ND2S U25023 ( .I1(n15888), .I2(n20359), .O(n19109) );
  ND2S U25024 ( .I1(n19110), .I2(n19109), .O(n13986) );
  MUX2S U25025 ( .A(n29587), .B(n20843), .S(gray_img[1312]), .O(n19112) );
  ND2S U25026 ( .I1(n15888), .I2(n20843), .O(n19111) );
  ND2S U25027 ( .I1(n19112), .I2(n19111), .O(n13998) );
  ND2S U25028 ( .I1(n15888), .I2(n20862), .O(n19113) );
  ND2S U25029 ( .I1(n19114), .I2(n19113), .O(n13853) );
  ND2S U25030 ( .I1(n15888), .I2(n20746), .O(n19115) );
  ND2S U25031 ( .I1(n19116), .I2(n19115), .O(n13826) );
  ND2S U25032 ( .I1(n15888), .I2(n20827), .O(n19117) );
  ND2S U25033 ( .I1(n19118), .I2(n19117), .O(n13894) );
  ND2S U25034 ( .I1(n15888), .I2(n20787), .O(n19119) );
  ND2S U25035 ( .I1(n19120), .I2(n19119), .O(n13895) );
  ND2S U25036 ( .I1(n15888), .I2(n20849), .O(n19121) );
  ND2S U25037 ( .I1(n19122), .I2(n19121), .O(n13827) );
  ND2S U25038 ( .I1(n15888), .I2(n20814), .O(n19123) );
  ND2S U25039 ( .I1(n19124), .I2(n19123), .O(n13967) );
  ND2S U25040 ( .I1(n15888), .I2(n20709), .O(n19125) );
  ND2S U25041 ( .I1(n19126), .I2(n19125), .O(n13958) );
  OA12S U25042 ( .B1(gray_img[423]), .B2(n29427), .A1(n27222), .O(n19129) );
  MOAI1S U25043 ( .A1(n27222), .A2(gray_img[423]), .B1(n25291), .B2(n19129), 
        .O(n19132) );
  NR2 U25044 ( .I1(gray_img[975]), .I2(gray_img[847]), .O(n23001) );
  INV1S U25045 ( .I(n23001), .O(n19130) );
  OR2S U25046 ( .I1(gray_img[839]), .I2(gray_img[967]), .O(n23000) );
  OAI12HS U25047 ( .B1(n19130), .B2(n23000), .A1(n15869), .O(n19131) );
  ND2S U25048 ( .I1(n19132), .I2(n19131), .O(n14118) );
  ND2S U25049 ( .I1(n15888), .I2(n20743), .O(n19133) );
  ND2S U25050 ( .I1(n19134), .I2(n19133), .O(n14082) );
  ND2S U25051 ( .I1(n15888), .I2(n20463), .O(n19135) );
  ND2S U25052 ( .I1(n19136), .I2(n19135), .O(n13910) );
  ND2S U25053 ( .I1(n15888), .I2(n20376), .O(n19137) );
  ND2S U25054 ( .I1(n19138), .I2(n19137), .O(n13859) );
  MUX2S U25055 ( .A(n30005), .B(n20559), .S(gray_img[880]), .O(n19140) );
  ND2S U25056 ( .I1(n15888), .I2(n20559), .O(n19139) );
  ND2S U25057 ( .I1(n19140), .I2(n19139), .O(n14128) );
  ND2S U25058 ( .I1(n15888), .I2(n20427), .O(n19141) );
  ND2S U25059 ( .I1(n19142), .I2(n19141), .O(n14001) );
  ND2S U25060 ( .I1(n15888), .I2(n20517), .O(n19143) );
  ND2S U25061 ( .I1(n19144), .I2(n19143), .O(n13988) );
  MUX2S U25062 ( .A(n30005), .B(n20562), .S(gray_img[1008]), .O(n19146) );
  ND2S U25063 ( .I1(n15888), .I2(n20562), .O(n19145) );
  ND2S U25064 ( .I1(n19146), .I2(n19145), .O(n14099) );
  MUX2S U25065 ( .A(n30050), .B(n20209), .S(gray_img[1984]), .O(n19148) );
  ND2S U25066 ( .I1(n15888), .I2(n20209), .O(n19147) );
  ND2S U25067 ( .I1(n19148), .I2(n19147), .O(n13823) );
  ND2S U25068 ( .I1(n15888), .I2(n20725), .O(n19149) );
  ND2S U25069 ( .I1(n19150), .I2(n19149), .O(n14011) );
  MUX2S U25070 ( .A(n30005), .B(n20365), .S(gray_img[744]), .O(n19152) );
  ND2S U25071 ( .I1(n15888), .I2(n20365), .O(n19151) );
  ND2S U25072 ( .I1(n19152), .I2(n19151), .O(n14151) );
  ND2S U25073 ( .I1(n15888), .I2(n20591), .O(n19153) );
  ND2S U25074 ( .I1(n19154), .I2(n19153), .O(n14178) );
  ND2S U25075 ( .I1(n15888), .I2(n20449), .O(n19155) );
  ND2S U25076 ( .I1(n19156), .I2(n19155), .O(n13870) );
  MUX2S U25077 ( .A(n30044), .B(n20602), .S(gray_img[1552]), .O(n19158) );
  ND2S U25078 ( .I1(n15888), .I2(n20602), .O(n19157) );
  ND2S U25079 ( .I1(n19158), .I2(n19157), .O(n13921) );
  ND2S U25080 ( .I1(n15888), .I2(n20550), .O(n19159) );
  ND2S U25081 ( .I1(n19160), .I2(n19159), .O(n13922) );
  ND2S U25082 ( .I1(n15888), .I2(n20440), .O(n19161) );
  ND2S U25083 ( .I1(n19162), .I2(n19161), .O(n13935) );
  MUX2S U25084 ( .A(n29032), .B(n20596), .S(gray_img[1560]), .O(n19164) );
  ND2S U25085 ( .I1(n15888), .I2(n20596), .O(n19163) );
  ND2S U25086 ( .I1(n19164), .I2(n19163), .O(n13920) );
  ND2S U25087 ( .I1(n15888), .I2(n20528), .O(n19165) );
  ND2S U25088 ( .I1(n19166), .I2(n19165), .O(n13915) );
  ND2S U25089 ( .I1(n15888), .I2(n20531), .O(n19167) );
  ND2S U25090 ( .I1(n19168), .I2(n19167), .O(n13906) );
  ND2S U25091 ( .I1(n15888), .I2(n20684), .O(n19169) );
  ND2S U25092 ( .I1(n19170), .I2(n19169), .O(n13951) );
  MUX2S U25093 ( .A(n20808), .B(n20054), .S(gray_img[752]), .O(n19172) );
  ND2S U25094 ( .I1(n15888), .I2(n20054), .O(n19171) );
  ND2S U25095 ( .I1(n19172), .I2(n19171), .O(n14143) );
  ND2S U25096 ( .I1(n15888), .I2(n25942), .O(n19174) );
  MUX2S U25097 ( .A(n30005), .B(n25942), .S(gray_img[2032]), .O(n19173) );
  ND2S U25098 ( .I1(n19174), .I2(n19173), .O(n13813) );
  ND2S U25099 ( .I1(n15888), .I2(n20509), .O(n19176) );
  ND2S U25100 ( .I1(n19176), .I2(n19175), .O(n13908) );
  MUX2S U25101 ( .A(n30005), .B(n20099), .S(gray_img[1020]), .O(n19177) );
  ND2S U25102 ( .I1(n19178), .I2(n19177), .O(n15005) );
  ND2S U25103 ( .I1(n19180), .I2(n19179), .O(n14987) );
  MUX2S U25104 ( .A(n20830), .B(n20512), .S(gray_img[1524]), .O(n19181) );
  ND2S U25105 ( .I1(n19184), .I2(n19183), .O(n14957) );
  MUX2S U25106 ( .A(n30005), .B(n20559), .S(gray_img[884]), .O(n19185) );
  ND2S U25107 ( .I1(n19186), .I2(n19185), .O(n15014) );
  MUX2S U25108 ( .A(n30005), .B(n20568), .S(gray_img[764]), .O(n19187) );
  ND2S U25109 ( .I1(n19188), .I2(n19187), .O(n15021) );
  MUX2S U25110 ( .A(n25928), .B(n20452), .S(gray_img[892]), .O(n19189) );
  ND2S U25111 ( .I1(n19190), .I2(n19189), .O(n15013) );
  MUX2S U25112 ( .A(n20808), .B(n20517), .S(gray_img[1396]), .O(n19191) );
  MUX2S U25113 ( .A(n20842), .B(n20035), .S(gray_img[1420]), .O(n19193) );
  MUX2S U25114 ( .A(n30005), .B(n20562), .S(gray_img[1012]), .O(n19195) );
  ND2S U25115 ( .I1(n19196), .I2(n19195), .O(n15006) );
  ND2S U25116 ( .I1(n19198), .I2(n19197), .O(n15061) );
  MUX2S U25117 ( .A(n20842), .B(n20427), .S(gray_img[1292]), .O(n19199) );
  MUX2S U25118 ( .A(n15904), .B(n20054), .S(gray_img[756]), .O(n19201) );
  ND2S U25119 ( .I1(n19202), .I2(n19201), .O(n15022) );
  ND2S U25120 ( .I1(n19204), .I2(n19203), .O(n14941) );
  ND2S U25121 ( .I1(n19206), .I2(n19205), .O(n14907) );
  MUX2S U25122 ( .A(n20808), .B(n20522), .S(gray_img[372]), .O(n19207) );
  ND2S U25123 ( .I1(n19208), .I2(n19207), .O(n15046) );
  ND2S U25124 ( .I1(n19210), .I2(n19209), .O(n14923) );
  MUX2S U25125 ( .A(n29587), .B(n20550), .S(gray_img[1548]), .O(n19211) );
  ND2S U25126 ( .I1(n19212), .I2(n19211), .O(n14939) );
  ND2S U25127 ( .I1(n19214), .I2(n19213), .O(n14926) );
  ND2S U25128 ( .I1(n19216), .I2(n19215), .O(n14900) );
  ND2S U25129 ( .I1(n19218), .I2(n19217), .O(n14895) );
  ND2S U25130 ( .I1(n19220), .I2(n19219), .O(n14932) );
  MUX2S U25131 ( .A(n30005), .B(n20463), .S(gray_img[1644]), .O(n19221) );
  ND2S U25132 ( .I1(n19222), .I2(n19221), .O(n14927) );
  MUX2S U25133 ( .A(n15904), .B(n20486), .S(gray_img[380]), .O(n19223) );
  ND2S U25134 ( .I1(n19224), .I2(n19223), .O(n15045) );
  MUX2S U25135 ( .A(n29032), .B(n20509), .S(gray_img[1660]), .O(n19225) );
  ND2S U25136 ( .I1(n19226), .I2(n19225), .O(n14925) );
  ND2S U25137 ( .I1(n19228), .I2(n19227), .O(n14893) );
  ND2S U25138 ( .I1(n19230), .I2(n19229), .O(n14891) );
  ND2S U25139 ( .I1(n19232), .I2(n19231), .O(n14909) );
  ND2S U25140 ( .I1(n19234), .I2(n19233), .O(n14916) );
  ND2S U25141 ( .I1(n19236), .I2(n19235), .O(n15030) );
  ND2S U25142 ( .I1(n19238), .I2(n19237), .O(n14910) );
  MUX2S U25143 ( .A(n25928), .B(n20565), .S(gray_img[636]), .O(n19239) );
  ND2S U25144 ( .I1(n19240), .I2(n19239), .O(n15029) );
  ND2S U25145 ( .I1(n19242), .I2(n19241), .O(n15037) );
  ND2S U25146 ( .I1(n19244), .I2(n19243), .O(n15053) );
  ND2S U25147 ( .I1(n19246), .I2(n19245), .O(n14911) );
  MUX2S U25148 ( .A(n29032), .B(n20063), .S(gray_img[1908]), .O(n19247) );
  ND2S U25149 ( .I1(n19248), .I2(n19247), .O(n14894) );
  MUX2S U25150 ( .A(n20842), .B(n20477), .S(gray_img[500]), .O(n19249) );
  MUX2S U25151 ( .A(n30005), .B(n20365), .S(gray_img[748]), .O(n19262) );
  MUX2S U25152 ( .A(n29566), .B(n20209), .S(gray_img[1988]), .O(n19264) );
  MUX2S U25153 ( .A(n30005), .B(n20142), .S(gray_img[1836]), .O(n19268) );
  MUX2S U25154 ( .A(n30005), .B(n20202), .S(gray_img[1964]), .O(n19270) );
  MUX2S U25155 ( .A(n30005), .B(n20212), .S(gray_img[876]), .O(n19272) );
  MUX2S U25156 ( .A(n30005), .B(n20129), .S(gray_img[1308]), .O(n19274) );
  MUX2S U25157 ( .A(n30005), .B(n20156), .S(gray_img[1828]), .O(n19276) );
  MUX2S U25158 ( .A(n30005), .B(n20384), .S(gray_img[1004]), .O(n19306) );
  MUX2S U25159 ( .A(n30005), .B(n20147), .S(gray_img[324]), .O(n19308) );
  ND2S U25160 ( .I1(n15888), .I2(n20857), .O(n19311) );
  ND2S U25161 ( .I1(n19312), .I2(n19311), .O(n14047) );
  ND2S U25162 ( .I1(n15888), .I2(n20193), .O(n19313) );
  ND2S U25163 ( .I1(n19314), .I2(n19313), .O(n13977) );
  ND2S U25164 ( .I1(n15888), .I2(n20395), .O(n19315) );
  ND2S U25165 ( .I1(n19316), .I2(n19315), .O(n13918) );
  ND2S U25166 ( .I1(n15888), .I2(n20392), .O(n19317) );
  ND2S U25167 ( .I1(n19318), .I2(n19317), .O(n14002) );
  MUX2S U25168 ( .A(n30050), .B(n20811), .S(gray_img[1440]), .O(n19320) );
  ND2S U25169 ( .I1(n15888), .I2(n20811), .O(n19319) );
  ND2S U25170 ( .I1(n19320), .I2(n19319), .O(n13968) );
  ND2S U25171 ( .I1(n15888), .I2(n20824), .O(n19321) );
  ND2S U25172 ( .I1(n19322), .I2(n19321), .O(n13919) );
  ND2S U25173 ( .I1(n15888), .I2(n20035), .O(n19323) );
  ND2S U25174 ( .I1(n19324), .I2(n19323), .O(n13985) );
  ND2S U25175 ( .I1(n15888), .I2(n20731), .O(n19325) );
  ND2S U25176 ( .I1(n19326), .I2(n19325), .O(n13916) );
  ND2S U25177 ( .I1(n15888), .I2(n20846), .O(n19327) );
  ND2S U25178 ( .I1(n19328), .I2(n19327), .O(n13889) );
  MUX2S U25179 ( .A(n30005), .B(n20129), .S(gray_img[1304]), .O(n19330) );
  ND2S U25180 ( .I1(n15888), .I2(n20129), .O(n19329) );
  ND2S U25181 ( .I1(n19330), .I2(n19329), .O(n13999) );
  MUX2S U25182 ( .A(n30005), .B(n20605), .S(gray_img[1680]), .O(n19332) );
  ND2S U25183 ( .I1(n15888), .I2(n20605), .O(n19331) );
  ND2S U25184 ( .I1(n19332), .I2(n19331), .O(n13901) );
  ND2S U25185 ( .I1(n15888), .I2(n20424), .O(n19333) );
  ND2S U25186 ( .I1(n19334), .I2(n19333), .O(n13842) );
  ND2S U25187 ( .I1(n15888), .I2(n20740), .O(n19335) );
  ND2S U25188 ( .I1(n19336), .I2(n19335), .O(n13852) );
  ND2S U25189 ( .I1(n15888), .I2(n20296), .O(n19337) );
  ND2S U25190 ( .I1(n19338), .I2(n19337), .O(n13856) );
  ND2S U25191 ( .I1(n15888), .I2(n20389), .O(n19339) );
  ND2S U25192 ( .I1(n19340), .I2(n19339), .O(n13837) );
  ND2S U25193 ( .I1(n15888), .I2(n20319), .O(n19341) );
  ND2S U25194 ( .I1(n19342), .I2(n19341), .O(n13858) );
  ND2S U25195 ( .I1(n15888), .I2(n19970), .O(n19343) );
  ND2S U25196 ( .I1(n19344), .I2(n19343), .O(n13836) );
  ND2S U25197 ( .I1(n15888), .I2(n20836), .O(n19345) );
  ND2S U25198 ( .I1(n19346), .I2(n19345), .O(n13997) );
  ND2S U25199 ( .I1(n19348), .I2(n19347), .O(n14948) );
  ND2S U25200 ( .I1(n19350), .I2(n19349), .O(n14996) );
  ND2S U25201 ( .I1(n19352), .I2(n19351), .O(n14885) );
  ND2S U25202 ( .I1(n19354), .I2(n19353), .O(n14959) );
  ND2S U25203 ( .I1(n19356), .I2(n19355), .O(n14917) );
  ND2S U25204 ( .I1(n19358), .I2(n19357), .O(n14933) );
  ND2S U25205 ( .I1(n19360), .I2(n19359), .O(n14975) );
  ND2S U25206 ( .I1(n19362), .I2(n19361), .O(n14973) );
  ND2S U25207 ( .I1(n19364), .I2(n19363), .O(n14991) );
  ND2S U25208 ( .I1(n19366), .I2(n19365), .O(n14989) );
  ND2S U25209 ( .I1(n19368), .I2(n19367), .O(n14901) );
  ND2S U25210 ( .I1(n19370), .I2(n19369), .O(n14943) );
  ND2S U25211 ( .I1(n19372), .I2(n19371), .O(n14918) );
  ND2S U25212 ( .I1(n19374), .I2(n19373), .O(n14935) );
  MUX2S U25213 ( .A(n15904), .B(n20811), .S(gray_img[1444]), .O(n19376) );
  ND2S U25214 ( .I1(n19376), .I2(n19375), .O(n14952) );
  ND2S U25215 ( .I1(n19378), .I2(n19377), .O(n14902) );
  ND2S U25216 ( .I1(n19380), .I2(n19379), .O(n14920) );
  ND2S U25217 ( .I1(n19382), .I2(n19381), .O(n14951) );
  ND2S U25218 ( .I1(n19384), .I2(n19383), .O(n14936) );
  ND2S U25219 ( .I1(n19386), .I2(n19385), .O(n14968) );
  ND2S U25220 ( .I1(n19388), .I2(n19387), .O(n14934) );
  ND2S U25221 ( .I1(n19390), .I2(n19389), .O(n14919) );
  ND2S U25222 ( .I1(n19392), .I2(n19391), .O(n14967) );
  ND2S U25223 ( .I1(n19394), .I2(n19393), .O(n14886) );
  OR2S U25224 ( .I1(n19396), .I2(n19402), .O(n19395) );
  NR2 U25225 ( .I1(n19395), .I2(n19403), .O(n24955) );
  INV1S U25226 ( .I(n19396), .O(n19401) );
  INV1S U25227 ( .I(n19397), .O(n19398) );
  NR2 U25228 ( .I1(n19398), .I2(n24944), .O(n24945) );
  OAI12HS U25229 ( .B1(n19401), .B2(n30360), .A1(n24949), .O(n24952) );
  NR2 U25230 ( .I1(n24955), .I2(n24952), .O(n25035) );
  INV1S U25231 ( .I(n25035), .O(n19399) );
  ND2S U25232 ( .I1(n19399), .I2(cnt_cro_y[0]), .O(n19405) );
  NR2 U25233 ( .I1(n19404), .I2(n19403), .O(n25041) );
  INV1S U25234 ( .I(cnt_cro_y[0]), .O(n30373) );
  ND2S U25235 ( .I1(n19405), .I2(n25034), .O(n15748) );
  AOI22S U25236 ( .A1(n19788), .A2(n19407), .B1(n25061), .B2(n19406), .O(
        n19408) );
  MUX2S U25237 ( .A(n30005), .B(n20614), .S(gray_img[2044]), .O(n19409) );
  ND2S U25238 ( .I1(n19410), .I2(n19409), .O(n14877) );
  ND2S U25239 ( .I1(n26828), .I2(n20614), .O(n19412) );
  MUX2S U25240 ( .A(n30005), .B(n20614), .S(gray_img[2045]), .O(n19411) );
  ND2S U25241 ( .I1(n19412), .I2(n19411), .O(n15077) );
  ND2S U25242 ( .I1(n15888), .I2(n20614), .O(n19414) );
  MUX2S U25243 ( .A(n30005), .B(n20614), .S(gray_img[2040]), .O(n19413) );
  ND2S U25244 ( .I1(n19414), .I2(n19413), .O(n13812) );
  AOI22S U25245 ( .A1(n25326), .A2(n19772), .B1(n25325), .B2(n25300), .O(
        n19415) );
  ND2S U25246 ( .I1(n25389), .I2(n20235), .O(n19417) );
  ND2S U25247 ( .I1(n19417), .I2(n19416), .O(n15399) );
  ND2S U25248 ( .I1(n26828), .I2(n20235), .O(n19419) );
  ND2S U25249 ( .I1(n19419), .I2(n19418), .O(n15203) );
  ND2S U25250 ( .I1(n19421), .I2(n19420), .O(n15003) );
  ND2S U25251 ( .I1(n19423), .I2(n19422), .O(n14403) );
  ND2S U25252 ( .I1(n15888), .I2(n20235), .O(n19425) );
  ND2S U25253 ( .I1(n19425), .I2(n19424), .O(n14089) );
  ND2S U25254 ( .I1(n15882), .I2(n20553), .O(n19427) );
  ND2S U25255 ( .I1(n19427), .I2(n19426), .O(n14588) );
  ND2S U25256 ( .I1(n15882), .I2(n20099), .O(n19429) );
  ND2S U25257 ( .I1(n19429), .I2(n19428), .O(n14606) );
  ND2S U25258 ( .I1(n15882), .I2(n20568), .O(n19431) );
  ND2S U25259 ( .I1(n19431), .I2(n19430), .O(n14622) );
  ND2S U25260 ( .I1(n15882), .I2(n20054), .O(n19433) );
  ND2S U25261 ( .I1(n19433), .I2(n19432), .O(n14623) );
  ND2S U25262 ( .I1(n15882), .I2(n20565), .O(n19435) );
  ND2S U25263 ( .I1(n19435), .I2(n19434), .O(n14630) );
  ND2S U25264 ( .I1(n15882), .I2(n20517), .O(n19437) );
  MUX2S U25265 ( .A(n20830), .B(n20517), .S(gray_img[1394]), .O(n19436) );
  ND2S U25266 ( .I1(n19437), .I2(n19436), .O(n14559) );
  ND2S U25267 ( .I1(n15881), .I2(n20544), .O(n19439) );
  ND2S U25268 ( .I1(n19439), .I2(n19438), .O(n14696) );
  ND2S U25269 ( .I1(n15882), .I2(n20571), .O(n19441) );
  ND2S U25270 ( .I1(n19441), .I2(n19440), .O(n14558) );
  ND2S U25271 ( .I1(n15881), .I2(n20504), .O(n19443) );
  ND2S U25272 ( .I1(n19443), .I2(n19442), .O(n14701) );
  ND2S U25273 ( .I1(n15882), .I2(n20512), .O(n19445) );
  MUX2S U25274 ( .A(n30005), .B(n20512), .S(gray_img[1522]), .O(n19444) );
  ND2S U25275 ( .I1(n19445), .I2(n19444), .O(n14543) );
  ND2S U25276 ( .I1(n15939), .I2(n20556), .O(n19447) );
  ND2S U25277 ( .I1(n19447), .I2(n19446), .O(n14542) );
  ND2S U25278 ( .I1(n15939), .I2(n20528), .O(n19449) );
  ND2S U25279 ( .I1(n19449), .I2(n19448), .O(n14533) );
  ND2S U25280 ( .I1(n15881), .I2(n20319), .O(n19451) );
  ND2S U25281 ( .I1(n19451), .I2(n19450), .O(n14708) );
  ND2S U25282 ( .I1(n15939), .I2(n20463), .O(n19453) );
  ND2S U25283 ( .I1(n19453), .I2(n19452), .O(n14528) );
  ND2S U25284 ( .I1(n15939), .I2(n19955), .O(n19455) );
  ND2S U25285 ( .I1(n19455), .I2(n19454), .O(n14517) );
  ND2S U25286 ( .I1(n15881), .I2(n20449), .O(n19457) );
  ND2S U25287 ( .I1(n19457), .I2(n19456), .O(n14712) );
  ND2S U25288 ( .I1(n15939), .I2(n20449), .O(n19459) );
  ND2S U25289 ( .I1(n19459), .I2(n19458), .O(n14512) );
  ND2S U25290 ( .I1(n15939), .I2(n20319), .O(n19461) );
  ND2S U25291 ( .I1(n19461), .I2(n19460), .O(n14508) );
  ND2S U25292 ( .I1(n15884), .I2(n20082), .O(n19463) );
  ND2S U25293 ( .I1(n19463), .I2(n19462), .O(n14461) );
  ND2S U25294 ( .I1(n15880), .I2(n19955), .O(n19465) );
  ND2S U25295 ( .I1(n19465), .I2(n19464), .O(n14717) );
  ND2S U25296 ( .I1(n15881), .I2(n20463), .O(n19467) );
  ND2S U25297 ( .I1(n19467), .I2(n19466), .O(n14728) );
  ND2S U25298 ( .I1(n15939), .I2(n20504), .O(n19469) );
  ND2S U25299 ( .I1(n19469), .I2(n19468), .O(n14501) );
  ND2S U25300 ( .I1(n15939), .I2(n20544), .O(n19471) );
  ND2S U25301 ( .I1(n19471), .I2(n19470), .O(n14496) );
  ND2S U25302 ( .I1(n15939), .I2(n20063), .O(n19473) );
  MUX2S U25303 ( .A(n20830), .B(n20063), .S(gray_img[1906]), .O(n19472) );
  ND2S U25304 ( .I1(n19473), .I2(n19472), .O(n14495) );
  ND2S U25305 ( .I1(n15939), .I2(n20430), .O(n19475) );
  ND2S U25306 ( .I1(n19475), .I2(n19474), .O(n14494) );
  ND2S U25307 ( .I1(n15883), .I2(n20424), .O(n19477) );
  ND2S U25308 ( .I1(n19477), .I2(n19476), .O(n14492) );
  ND2S U25309 ( .I1(n15880), .I2(n20528), .O(n19479) );
  ND2S U25310 ( .I1(n19479), .I2(n19478), .O(n14733) );
  ND2S U25311 ( .I1(n15884), .I2(n20486), .O(n19481) );
  ND2S U25312 ( .I1(n19481), .I2(n19480), .O(n14445) );
  ND2S U25313 ( .I1(n15885), .I2(n20559), .O(n19483) );
  ND2S U25314 ( .I1(n19483), .I2(n19482), .O(n14414) );
  ND2S U25315 ( .I1(n15933), .I2(n20562), .O(n19485) );
  ND2S U25316 ( .I1(n19485), .I2(n19484), .O(n14406) );
  ND2S U25317 ( .I1(n15933), .I2(n20496), .O(n19487) );
  ND2S U25318 ( .I1(n19487), .I2(n19486), .O(n14453) );
  ND2S U25319 ( .I1(n15881), .I2(n20099), .O(n19489) );
  ND2S U25320 ( .I1(n19489), .I2(n19488), .O(n14806) );
  ND2S U25321 ( .I1(n15885), .I2(n20556), .O(n19491) );
  ND2S U25322 ( .I1(n19491), .I2(n19490), .O(n14341) );
  ND2S U25323 ( .I1(n15933), .I2(n20472), .O(n19493) );
  MUX2S U25324 ( .A(n20830), .B(n20472), .S(gray_img[505]), .O(n19492) );
  ND2S U25325 ( .I1(n19493), .I2(n19492), .O(n14437) );
  ND2S U25326 ( .I1(n15880), .I2(n20568), .O(n19495) );
  ND2S U25327 ( .I1(n19495), .I2(n19494), .O(n14822) );
  ND2S U25328 ( .I1(n15880), .I2(n20054), .O(n19497) );
  ND2S U25329 ( .I1(n19497), .I2(n19496), .O(n14823) );
  ND2S U25330 ( .I1(n15926), .I2(n20565), .O(n19499) );
  ND2S U25331 ( .I1(n19499), .I2(n19498), .O(n14830) );
  ND2S U25332 ( .I1(n15933), .I2(n20517), .O(n19501) );
  MUX2S U25333 ( .A(n20830), .B(n20517), .S(gray_img[1393]), .O(n19500) );
  ND2S U25334 ( .I1(n19501), .I2(n19500), .O(n14358) );
  ND2S U25335 ( .I1(n15933), .I2(n20571), .O(n19503) );
  ND2S U25336 ( .I1(n19503), .I2(n19502), .O(n14357) );
  ND2S U25337 ( .I1(n15933), .I2(n20553), .O(n19505) );
  ND2S U25338 ( .I1(n19505), .I2(n19504), .O(n14387) );
  ND2S U25339 ( .I1(n15880), .I2(n20472), .O(n19507) );
  MUX2S U25340 ( .A(n30005), .B(n20472), .S(gray_img[507]), .O(n19506) );
  ND2S U25341 ( .I1(n19507), .I2(n19506), .O(n14838) );
  ND2S U25342 ( .I1(n15880), .I2(n20477), .O(n19509) );
  ND2S U25343 ( .I1(n19509), .I2(n19508), .O(n14839) );
  ND2S U25344 ( .I1(n15881), .I2(n20486), .O(n19511) );
  ND2S U25345 ( .I1(n19511), .I2(n19510), .O(n14846) );
  ND2S U25346 ( .I1(n15881), .I2(n20496), .O(n19513) );
  ND2S U25347 ( .I1(n19513), .I2(n19512), .O(n14854) );
  ND2S U25348 ( .I1(n15933), .I2(n20512), .O(n19515) );
  ND2S U25349 ( .I1(n19515), .I2(n19514), .O(n14342) );
  ND2S U25350 ( .I1(n15933), .I2(n20550), .O(n19517) );
  ND2S U25351 ( .I1(n19517), .I2(n19516), .O(n14339) );
  ND2S U25352 ( .I1(n15933), .I2(n20099), .O(n19519) );
  ND2S U25353 ( .I1(n19519), .I2(n19518), .O(n14405) );
  ND2S U25354 ( .I1(n15884), .I2(n20452), .O(n19521) );
  ND2S U25355 ( .I1(n19521), .I2(n19520), .O(n14413) );
  ND2S U25356 ( .I1(n15880), .I2(n20082), .O(n19523) );
  ND2S U25357 ( .I1(n19523), .I2(n19522), .O(n14862) );
  ND2S U25358 ( .I1(n15880), .I2(n20424), .O(n19525) );
  ND2S U25359 ( .I1(n19525), .I2(n19524), .O(n14692) );
  ND2S U25360 ( .I1(n15884), .I2(n20477), .O(n19527) );
  ND2S U25361 ( .I1(n19527), .I2(n19526), .O(n14438) );
  ND2S U25362 ( .I1(n15928), .I2(n19955), .O(n19529) );
  ND2S U25363 ( .I1(n19529), .I2(n19528), .O(n14316) );
  ND2S U25364 ( .I1(n15928), .I2(n20054), .O(n19531) );
  ND2S U25365 ( .I1(n19531), .I2(n19530), .O(n14422) );
  ND2S U25366 ( .I1(n15885), .I2(n20534), .O(n19533) );
  ND2S U25367 ( .I1(n19533), .I2(n19532), .O(n14430) );
  ND2S U25368 ( .I1(n15884), .I2(n20463), .O(n19535) );
  ND2S U25369 ( .I1(n19535), .I2(n19534), .O(n14327) );
  ND2S U25370 ( .I1(n15885), .I2(n20449), .O(n19537) );
  ND2S U25371 ( .I1(n19537), .I2(n19536), .O(n14311) );
  ND2S U25372 ( .I1(n15884), .I2(n20531), .O(n19539) );
  ND2S U25373 ( .I1(n19539), .I2(n19538), .O(n14323) );
  ND2S U25374 ( .I1(n15880), .I2(n19970), .O(n19540) );
  ND2S U25375 ( .I1(n19541), .I2(n19540), .O(n14690) );
  ND2S U25376 ( .I1(n15884), .I2(n20596), .O(n19542) );
  ND2S U25377 ( .I1(n19543), .I2(n19542), .O(n14337) );
  MUX2S U25378 ( .A(n30005), .B(n20129), .S(gray_img[1307]), .O(n19545) );
  ND2S U25379 ( .I1(n15887), .I2(n20129), .O(n19544) );
  ND2S U25380 ( .I1(n19545), .I2(n19544), .O(n14770) );
  ND2S U25381 ( .I1(n15887), .I2(n20184), .O(n19546) );
  ND2S U25382 ( .I1(n19547), .I2(n19546), .O(n14802) );
  ND2S U25383 ( .I1(n15884), .I2(n20602), .O(n19548) );
  ND2S U25384 ( .I1(n19549), .I2(n19548), .O(n14338) );
  MUX2S U25385 ( .A(n30005), .B(n20202), .S(gray_img[1962]), .O(n19551) );
  ND2S U25386 ( .I1(n15937), .I2(n20202), .O(n19550) );
  ND2S U25387 ( .I1(n19551), .I2(n19550), .O(n14488) );
  ND2S U25388 ( .I1(n15883), .I2(n20379), .O(n19552) );
  ND2S U25389 ( .I1(n19553), .I2(n19552), .O(n14585) );
  MUX2S U25390 ( .A(n30005), .B(n20129), .S(gray_img[1306]), .O(n19555) );
  ND2S U25391 ( .I1(n15883), .I2(n20129), .O(n19554) );
  ND2S U25392 ( .I1(n19555), .I2(n19554), .O(n14570) );
  ND2S U25393 ( .I1(n15884), .I2(n20583), .O(n19556) );
  ND2S U25394 ( .I1(n19557), .I2(n19556), .O(n14324) );
  ND2S U25395 ( .I1(n15887), .I2(n20373), .O(n19558) );
  ND2S U25396 ( .I1(n19559), .I2(n19558), .O(n14693) );
  MUX2S U25397 ( .A(n30005), .B(n20202), .S(gray_img[1963]), .O(n19561) );
  ND2S U25398 ( .I1(n15887), .I2(n20202), .O(n19560) );
  ND2S U25399 ( .I1(n19561), .I2(n19560), .O(n14688) );
  MUX2S U25400 ( .A(n30005), .B(n20147), .S(gray_img[322]), .O(n19563) );
  ND2S U25401 ( .I1(n15883), .I2(n20147), .O(n19562) );
  ND2S U25402 ( .I1(n19563), .I2(n19562), .O(n14653) );
  MUX2S U25403 ( .A(n30005), .B(n20384), .S(gray_img[1003]), .O(n19565) );
  ND2S U25404 ( .I1(n15887), .I2(n20384), .O(n19564) );
  ND2S U25405 ( .I1(n19565), .I2(n19564), .O(n14808) );
  ND2S U25406 ( .I1(n15883), .I2(n20193), .O(n19566) );
  ND2S U25407 ( .I1(n19567), .I2(n19566), .O(n14555) );
  ND2S U25408 ( .I1(n15884), .I2(n20293), .O(n19568) );
  ND2S U25409 ( .I1(n19569), .I2(n19568), .O(n14353) );
  ND2S U25410 ( .I1(n15884), .I2(n20193), .O(n19570) );
  ND2S U25411 ( .I1(n19571), .I2(n19570), .O(n14354) );
  ND2S U25412 ( .I1(n15939), .I2(n20591), .O(n19572) );
  ND2S U25413 ( .I1(n19573), .I2(n19572), .O(n14637) );
  ND2S U25414 ( .I1(n15887), .I2(n20389), .O(n19574) );
  ND2S U25415 ( .I1(n19575), .I2(n19574), .O(n14691) );
  MUX2S U25416 ( .A(n30005), .B(n20365), .S(gray_img[747]), .O(n19577) );
  ND2S U25417 ( .I1(n15887), .I2(n20365), .O(n19576) );
  ND2S U25418 ( .I1(n19577), .I2(n19576), .O(n14824) );
  MUX2S U25419 ( .A(n30005), .B(n20599), .S(gray_img[1689]), .O(n19579) );
  ND2S U25420 ( .I1(n15884), .I2(n20599), .O(n19578) );
  ND2S U25421 ( .I1(n19579), .I2(n19578), .O(n14321) );
  ND2S U25422 ( .I1(n15883), .I2(n20362), .O(n19580) );
  ND2S U25423 ( .I1(n19581), .I2(n19580), .O(n14571) );
  ND2S U25424 ( .I1(n15881), .I2(n20362), .O(n19582) );
  ND2S U25425 ( .I1(n19583), .I2(n19582), .O(n14771) );
  MUX2S U25426 ( .A(n30005), .B(n20147), .S(gray_img[323]), .O(n19585) );
  ND2S U25427 ( .I1(n15881), .I2(n20147), .O(n19584) );
  ND2S U25428 ( .I1(n19585), .I2(n19584), .O(n14853) );
  ND2S U25429 ( .I1(n15881), .I2(n20376), .O(n19586) );
  ND2S U25430 ( .I1(n19587), .I2(n19586), .O(n14709) );
  ND2S U25431 ( .I1(n15880), .I2(n20193), .O(n19588) );
  ND2S U25432 ( .I1(n19589), .I2(n19588), .O(n14755) );
  ND2S U25433 ( .I1(n15883), .I2(n20296), .O(n19590) );
  ND2S U25434 ( .I1(n19591), .I2(n19590), .O(n14506) );
  ND2S U25435 ( .I1(n15932), .I2(n20362), .O(n19592) );
  ND2S U25436 ( .I1(n19593), .I2(n19592), .O(n14370) );
  ND2S U25437 ( .I1(n15884), .I2(n20142), .O(n19594) );
  ND2S U25438 ( .I1(n19595), .I2(n19594), .O(n14303) );
  ND2S U25439 ( .I1(n15883), .I2(n20580), .O(n19596) );
  ND2S U25440 ( .I1(n19597), .I2(n19596), .O(n14613) );
  ND2S U25441 ( .I1(n15927), .I2(n20296), .O(n19598) );
  ND2S U25442 ( .I1(n19599), .I2(n19598), .O(n14706) );
  MUX2S U25443 ( .A(n30005), .B(n20384), .S(gray_img[1002]), .O(n19601) );
  ND2S U25444 ( .I1(n15937), .I2(n20384), .O(n19600) );
  ND2S U25445 ( .I1(n19601), .I2(n19600), .O(n14608) );
  ND2S U25446 ( .I1(n15937), .I2(n20184), .O(n19602) );
  ND2S U25447 ( .I1(n19603), .I2(n19602), .O(n14602) );
  MUX2S U25448 ( .A(n29587), .B(n20368), .S(gray_img[1058]), .O(n19605) );
  ND2S U25449 ( .I1(n15937), .I2(n20368), .O(n19604) );
  ND2S U25450 ( .I1(n19605), .I2(n19604), .O(n14601) );
  MUX2S U25451 ( .A(n30005), .B(n20147), .S(gray_img[321]), .O(n19607) );
  ND2S U25452 ( .I1(n15886), .I2(n20147), .O(n19606) );
  ND2S U25453 ( .I1(n19607), .I2(n19606), .O(n14452) );
  MUX2S U25454 ( .A(n30005), .B(n20373), .S(gray_img[1922]), .O(n19609) );
  ND2S U25455 ( .I1(n15937), .I2(n20373), .O(n19608) );
  ND2S U25456 ( .I1(n19609), .I2(n19608), .O(n14493) );
  ND2S U25457 ( .I1(n15886), .I2(n20184), .O(n19610) );
  ND2S U25458 ( .I1(n19611), .I2(n19610), .O(n14401) );
  MUX2S U25459 ( .A(n29032), .B(n20376), .S(gray_img[1794]), .O(n19613) );
  ND2S U25460 ( .I1(n15937), .I2(n20376), .O(n19612) );
  ND2S U25461 ( .I1(n19613), .I2(n19612), .O(n14509) );
  ND2S U25462 ( .I1(n15937), .I2(n19970), .O(n19614) );
  ND2S U25463 ( .I1(n19615), .I2(n19614), .O(n14490) );
  ND2S U25464 ( .I1(n15886), .I2(n20605), .O(n19616) );
  ND2S U25465 ( .I1(n19617), .I2(n19616), .O(n14322) );
  ND2S U25466 ( .I1(n15886), .I2(n20296), .O(n19618) );
  ND2S U25467 ( .I1(n19619), .I2(n19618), .O(n14305) );
  MUX2S U25468 ( .A(n30005), .B(n20156), .S(gray_img[1825]), .O(n19621) );
  ND2S U25469 ( .I1(n15931), .I2(n20156), .O(n19620) );
  ND2S U25470 ( .I1(n19621), .I2(n19620), .O(n14304) );
  MUX2S U25471 ( .A(n30005), .B(n20212), .S(gray_img[875]), .O(n19623) );
  ND2S U25472 ( .I1(n15927), .I2(n20212), .O(n19622) );
  ND2S U25473 ( .I1(n19623), .I2(n19622), .O(n14816) );
  MUX2S U25474 ( .A(n30005), .B(n20212), .S(gray_img[874]), .O(n19625) );
  ND2S U25475 ( .I1(n15937), .I2(n20212), .O(n19624) );
  ND2S U25476 ( .I1(n19625), .I2(n19624), .O(n14616) );
  ND2S U25477 ( .I1(n15937), .I2(n20389), .O(n19626) );
  ND2S U25478 ( .I1(n19627), .I2(n19626), .O(n14491) );
  MUX2S U25479 ( .A(n30005), .B(n20156), .S(gray_img[1826]), .O(n19629) );
  ND2S U25480 ( .I1(n15939), .I2(n20156), .O(n19628) );
  ND2S U25481 ( .I1(n19629), .I2(n19628), .O(n14505) );
  ND2S U25482 ( .I1(n15937), .I2(n25942), .O(n19631) );
  MUX2S U25483 ( .A(n30005), .B(n25942), .S(gray_img[2034]), .O(n19630) );
  ND2S U25484 ( .I1(n19631), .I2(n19630), .O(n14479) );
  ND2S U25485 ( .I1(n19633), .I2(n19632), .O(n14791) );
  ND2S U25486 ( .I1(n19635), .I2(n19634), .O(n14390) );
  ND2S U25487 ( .I1(n19637), .I2(n19636), .O(n14744) );
  ND2S U25488 ( .I1(n19639), .I2(n19638), .O(n14544) );
  ND2S U25489 ( .I1(n19641), .I2(n19640), .O(n14591) );
  ND2S U25490 ( .I1(n19643), .I2(n19642), .O(n14343) );
  ND2S U25491 ( .I1(n15927), .I2(n20235), .O(n19645) );
  ND2S U25492 ( .I1(n19645), .I2(n19644), .O(n14804) );
  ND2S U25493 ( .I1(n15937), .I2(n20614), .O(n19647) );
  MUX2S U25494 ( .A(n30005), .B(n20614), .S(gray_img[2042]), .O(n19646) );
  ND2S U25495 ( .I1(n19647), .I2(n19646), .O(n14478) );
  ND2S U25496 ( .I1(n15939), .I2(n20235), .O(n19649) );
  ND2S U25497 ( .I1(n19649), .I2(n19648), .O(n14604) );
  ND2S U25498 ( .I1(n15880), .I2(n20614), .O(n19651) );
  MUX2S U25499 ( .A(n30005), .B(n20614), .S(gray_img[2043]), .O(n19650) );
  ND2S U25500 ( .I1(n19651), .I2(n19650), .O(n14678) );
  ND2S U25501 ( .I1(n19653), .I2(n19652), .O(n14336) );
  ND2S U25502 ( .I1(n19655), .I2(n19654), .O(n14335) );
  ND2S U25503 ( .I1(n19657), .I2(n19656), .O(n14721) );
  ND2S U25504 ( .I1(n19659), .I2(n19658), .O(n14521) );
  ND2S U25505 ( .I1(n19661), .I2(n19660), .O(n14536) );
  ND2S U25506 ( .I1(n19663), .I2(n19662), .O(n14736) );
  AOI22S U25507 ( .A1(n25245), .A2(n19772), .B1(n25244), .B2(n25300), .O(
        n19664) );
  ND2S U25508 ( .I1(n15891), .I2(n20611), .O(n19666) );
  ND2S U25509 ( .I1(n19666), .I2(n19665), .O(n15199) );
  AOI22S U25510 ( .A1(n25245), .A2(n19758), .B1(n25244), .B2(n25296), .O(
        n19667) );
  ND2S U25511 ( .I1(n19669), .I2(n19668), .O(n14983) );
  ND2S U25512 ( .I1(n15891), .I2(n20435), .O(n19671) );
  ND2S U25513 ( .I1(n19671), .I2(n19670), .O(n15183) );
  ND2S U25514 ( .I1(n19673), .I2(n19672), .O(n14999) );
  ND2S U25515 ( .I1(n15888), .I2(n20435), .O(n19675) );
  ND2S U25516 ( .I1(n19675), .I2(n19674), .O(n14055) );
  ND2S U25517 ( .I1(n15888), .I2(n20611), .O(n19677) );
  ND2S U25518 ( .I1(n19677), .I2(n19676), .O(n14085) );
  ND2S U25519 ( .I1(n19679), .I2(n19678), .O(n14784) );
  ND2S U25520 ( .I1(n19681), .I2(n19680), .O(n14383) );
  ND2S U25521 ( .I1(n19683), .I2(n19682), .O(n14800) );
  ND2S U25522 ( .I1(n19685), .I2(n19684), .O(n14584) );
  ND2S U25523 ( .I1(n19687), .I2(n19686), .O(n14399) );
  AOI22S U25524 ( .A1(n25218), .A2(n19772), .B1(n25216), .B2(n25300), .O(
        n19688) );
  ND2S U25525 ( .I1(n26828), .I2(n20311), .O(n19690) );
  MUX2S U25526 ( .A(n30005), .B(n20311), .S(gray_img[1029]), .O(n19689) );
  ND2S U25527 ( .I1(n19690), .I2(n19689), .O(n15204) );
  ND2S U25528 ( .I1(n15884), .I2(n20311), .O(n19692) );
  MUX2S U25529 ( .A(n30005), .B(n20311), .S(gray_img[1025]), .O(n19691) );
  ND2S U25530 ( .I1(n19692), .I2(n19691), .O(n14404) );
  ND2S U25531 ( .I1(n15937), .I2(n20311), .O(n19694) );
  MUX2S U25532 ( .A(n30005), .B(n20311), .S(gray_img[1026]), .O(n19693) );
  ND2S U25533 ( .I1(n19694), .I2(n19693), .O(n14605) );
  ND2S U25534 ( .I1(n15927), .I2(n20311), .O(n19696) );
  MUX2S U25535 ( .A(n30005), .B(n20311), .S(gray_img[1027]), .O(n19695) );
  ND2S U25536 ( .I1(n19696), .I2(n19695), .O(n14805) );
  MUX2S U25537 ( .A(n30005), .B(n20311), .S(gray_img[1028]), .O(n19697) );
  ND2S U25538 ( .I1(n19698), .I2(n19697), .O(n15004) );
  AOI22S U25539 ( .A1(n25218), .A2(n19758), .B1(n25216), .B2(n25296), .O(
        n19699) );
  ND2S U25540 ( .I1(n15937), .I2(n20240), .O(n19701) );
  ND2S U25541 ( .I1(n19701), .I2(n19700), .O(n14589) );
  ND2S U25542 ( .I1(n26828), .I2(n20240), .O(n19703) );
  ND2S U25543 ( .I1(n19703), .I2(n19702), .O(n15188) );
  ND2S U25544 ( .I1(n19705), .I2(n19704), .O(n14988) );
  ND2S U25545 ( .I1(n15927), .I2(n20240), .O(n19707) );
  ND2S U25546 ( .I1(n19707), .I2(n19706), .O(n14789) );
  ND2S U25547 ( .I1(n15888), .I2(n20240), .O(n19709) );
  ND2S U25548 ( .I1(n19709), .I2(n19708), .O(n14074) );
  ND2S U25549 ( .I1(n15888), .I2(n20311), .O(n19711) );
  MUX2S U25550 ( .A(n30005), .B(n20311), .S(gray_img[1024]), .O(n19710) );
  ND2S U25551 ( .I1(n19711), .I2(n19710), .O(n14090) );
  ND2S U25552 ( .I1(n19713), .I2(n19712), .O(n14388) );
  AOI22S U25553 ( .A1(n25246), .A2(n19720), .B1(n25257), .B2(n19719), .O(
        n19714) );
  ND2S U25554 ( .I1(n15886), .I2(n20260), .O(n19716) );
  AOI22S U25555 ( .A1(n25273), .A2(n19720), .B1(n25271), .B2(n19719), .O(
        n19721) );
  ND2S U25556 ( .I1(n15891), .I2(n20499), .O(n19725) );
  AOI22S U25557 ( .A1(n25283), .A2(n19772), .B1(n25282), .B2(n25300), .O(
        n19726) );
  ND2S U25558 ( .I1(n15884), .I2(n20499), .O(n19730) );
  AOI22S U25559 ( .A1(n25283), .A2(n19758), .B1(n25282), .B2(n25296), .O(
        n19731) );
  ND2S U25560 ( .I1(n15890), .I2(n20260), .O(n19735) );
  ND2S U25561 ( .I1(n26828), .I2(n20260), .O(n19737) );
  ND2S U25562 ( .I1(n15888), .I2(n20757), .O(n19739) );
  ND2S U25563 ( .I1(n15891), .I2(n20757), .O(n19741) );
  ND2S U25564 ( .I1(n15891), .I2(n20760), .O(n19743) );
  ND2S U25565 ( .I1(n15888), .I2(n20760), .O(n19745) );
  ND2S U25566 ( .I1(n15888), .I2(n20260), .O(n19747) );
  ND2S U25567 ( .I1(n15888), .I2(n20499), .O(n19755) );
  MUX2S U25568 ( .A(n20842), .B(n20499), .S(gray_img[112]), .O(n19754) );
  AOI22S U25569 ( .A1(n25274), .A2(n19758), .B1(n25272), .B2(n25296), .O(
        n19759) );
  ND2S U25570 ( .I1(n26828), .I2(n20316), .O(n19761) );
  ND2S U25571 ( .I1(n19761), .I2(n19760), .O(n15186) );
  ND2S U25572 ( .I1(n19763), .I2(n19762), .O(n14986) );
  ND2S U25573 ( .I1(n15888), .I2(n20316), .O(n19765) );
  ND2S U25574 ( .I1(n19765), .I2(n19764), .O(n14065) );
  ND2S U25575 ( .I1(n19767), .I2(n19766), .O(n14386) );
  ND2S U25576 ( .I1(n19769), .I2(n19768), .O(n14587) );
  ND2S U25577 ( .I1(n19771), .I2(n19770), .O(n14787) );
  AOI22S U25578 ( .A1(n25274), .A2(n19772), .B1(n25272), .B2(n25300), .O(
        n19773) );
  ND2S U25579 ( .I1(n26445), .I2(n20255), .O(n19777) );
  ND2S U25580 ( .I1(n25389), .I2(n20255), .O(n19779) );
  ND2S U25581 ( .I1(n15888), .I2(n20255), .O(n19781) );
  AOI22S U25582 ( .A1(n19788), .A2(n19845), .B1(n25061), .B2(n19844), .O(
        n19789) );
  ND2S U25583 ( .I1(n15891), .I2(n20608), .O(n19791) );
  MUX2S U25584 ( .A(n30005), .B(n20608), .S(gray_img[2029]), .O(n19790) );
  ND2S U25585 ( .I1(n19791), .I2(n19790), .O(n15079) );
  ND2S U25586 ( .I1(n15937), .I2(n20608), .O(n19793) );
  MUX2S U25587 ( .A(n30005), .B(n20608), .S(gray_img[2026]), .O(n19792) );
  ND2S U25588 ( .I1(n19793), .I2(n19792), .O(n14480) );
  MUX2S U25589 ( .A(n30005), .B(n20608), .S(gray_img[2028]), .O(n19794) );
  ND2S U25590 ( .I1(n19795), .I2(n19794), .O(n14879) );
  ND2S U25591 ( .I1(n15880), .I2(n20608), .O(n19797) );
  MUX2S U25592 ( .A(n30005), .B(n20608), .S(gray_img[2027]), .O(n19796) );
  ND2S U25593 ( .I1(n19797), .I2(n19796), .O(n14680) );
  ND2S U25594 ( .I1(n15888), .I2(n20608), .O(n19799) );
  MUX2S U25595 ( .A(n30005), .B(n20608), .S(gray_img[2024]), .O(n19798) );
  ND2S U25596 ( .I1(n19799), .I2(n19798), .O(n13815) );
  AOI22S U25597 ( .A1(n25162), .A2(n19845), .B1(n25361), .B2(n19844), .O(
        n19800) );
  ND2S U25598 ( .I1(n27751), .I2(n20491), .O(n19802) );
  ND2S U25599 ( .I1(n19802), .I2(n19801), .O(n15247) );
  ND2S U25600 ( .I1(n19804), .I2(n19803), .O(n15047) );
  ND2S U25601 ( .I1(n15886), .I2(n20491), .O(n19806) );
  ND2S U25602 ( .I1(n19806), .I2(n19805), .O(n14447) );
  AOI22S U25603 ( .A1(n25372), .A2(n19845), .B1(n25370), .B2(n19844), .O(
        n19807) );
  ND2S U25604 ( .I1(n15931), .I2(n20480), .O(n19809) );
  ND2S U25605 ( .I1(n19809), .I2(n19808), .O(n14439) );
  ND2S U25606 ( .I1(n19811), .I2(n19810), .O(n15039) );
  ND2S U25607 ( .I1(n15891), .I2(n20480), .O(n19813) );
  ND2S U25608 ( .I1(n19813), .I2(n19812), .O(n15239) );
  ND2S U25609 ( .I1(n15888), .I2(n20491), .O(n19815) );
  ND2S U25610 ( .I1(n19815), .I2(n19814), .O(n14217) );
  ND2S U25611 ( .I1(n19817), .I2(n19816), .O(n14848) );
  ND2S U25612 ( .I1(n19819), .I2(n19818), .O(n14648) );
  ND2S U25613 ( .I1(n19821), .I2(n19820), .O(n14840) );
  ND2S U25614 ( .I1(n19823), .I2(n19822), .O(n14640) );
  ND2S U25615 ( .I1(n15888), .I2(n20480), .O(n19825) );
  ND2S U25616 ( .I1(n19825), .I2(n19824), .O(n14195) );
  AOI22S U25617 ( .A1(n25246), .A2(n19845), .B1(n25257), .B2(n19844), .O(
        n19826) );
  ND2S U25618 ( .I1(n15891), .I2(n20620), .O(n19828) );
  INV1S U25619 ( .I(gray_img[237]), .O(n27400) );
  MUX2S U25620 ( .A(n20620), .B(n30050), .S(n27400), .O(n19827) );
  ND2S U25621 ( .I1(n19828), .I2(n19827), .O(n15255) );
  ND2S U25622 ( .I1(n19830), .I2(n19829), .O(n15055) );
  ND2S U25623 ( .I1(n15881), .I2(n20620), .O(n19832) );
  ND2S U25624 ( .I1(n19832), .I2(n19831), .O(n14856) );
  AOI22S U25625 ( .A1(n25195), .A2(n19845), .B1(n25333), .B2(n19844), .O(
        n19833) );
  ND2S U25626 ( .I1(n15885), .I2(n20274), .O(n19837) );
  ND2S U25627 ( .I1(n15891), .I2(n20274), .O(n19839) );
  MUX2S U25628 ( .A(n30005), .B(n20274), .S(gray_img[621]), .O(n19838) );
  ND2S U25629 ( .I1(n25389), .I2(n20274), .O(n19841) );
  ND2S U25630 ( .I1(n19843), .I2(n19842), .O(n14656) );
  AOI22S U25631 ( .A1(n25273), .A2(n19845), .B1(n25271), .B2(n19844), .O(
        n19846) );
  ND2S U25632 ( .I1(n15891), .I2(n20617), .O(n19848) );
  INV1S U25633 ( .I(gray_img[109]), .O(n27402) );
  ND2S U25634 ( .I1(n19848), .I2(n19847), .O(n15263) );
  ND2S U25635 ( .I1(n15888), .I2(n20620), .O(n19854) );
  ND2S U25636 ( .I1(n19854), .I2(n19853), .O(n14239) );
  ND2S U25637 ( .I1(n15881), .I2(n20617), .O(n19856) );
  ND2S U25638 ( .I1(n19856), .I2(n19855), .O(n14864) );
  ND2S U25639 ( .I1(n19858), .I2(n19857), .O(n15063) );
  ND2S U25640 ( .I1(n15888), .I2(n20274), .O(n19860) );
  ND2S U25641 ( .I1(n19862), .I2(n19861), .O(n14664) );
  ND2S U25642 ( .I1(n15888), .I2(n20617), .O(n19864) );
  ND2S U25643 ( .I1(n19864), .I2(n19863), .O(n14261) );
  AOI22S U25644 ( .A1(n25308), .A2(n19914), .B1(n25340), .B2(n19913), .O(
        n19865) );
  ND2S U25645 ( .I1(n27751), .I2(n20623), .O(n19867) );
  ND2S U25646 ( .I1(n15887), .I2(n20623), .O(n19869) );
  ND2S U25647 ( .I1(n25389), .I2(n20623), .O(n19873) );
  AOI22S U25648 ( .A1(n25372), .A2(n19914), .B1(n25370), .B2(n19913), .O(
        n19874) );
  ND2S U25649 ( .I1(n15891), .I2(n20483), .O(n19876) );
  MUX2S U25650 ( .A(n25928), .B(n20483), .S(gray_img[453]), .O(n19875) );
  MUX2S U25651 ( .A(n25928), .B(n20483), .S(gray_img[452]), .O(n19877) );
  ND2S U25652 ( .I1(n15888), .I2(n20623), .O(n19880) );
  MUX2S U25653 ( .A(n25928), .B(n20623), .S(gray_img[706]), .O(n19881) );
  MUX2S U25654 ( .A(n25928), .B(n20483), .S(gray_img[449]), .O(n19883) );
  ND2S U25655 ( .I1(n15888), .I2(n20483), .O(n19886) );
  MUX2S U25656 ( .A(n25928), .B(n20483), .S(gray_img[448]), .O(n19885) );
  MUX2S U25657 ( .A(n25928), .B(n20483), .S(gray_img[451]), .O(n19887) );
  MUX2S U25658 ( .A(n25928), .B(n20483), .S(gray_img[450]), .O(n19889) );
  AOI22S U25659 ( .A1(n25246), .A2(n19914), .B1(n25257), .B2(n19913), .O(
        n19891) );
  ND2S U25660 ( .I1(n25389), .I2(n20631), .O(n19893) );
  ND2S U25661 ( .I1(n15880), .I2(n20631), .O(n19897) );
  ND2S U25662 ( .I1(n15891), .I2(n20631), .O(n19899) );
  ND2S U25663 ( .I1(n15888), .I2(n20631), .O(n19901) );
  AOI22S U25664 ( .A1(n25273), .A2(n19914), .B1(n25271), .B2(n19913), .O(
        n19904) );
  ND2S U25665 ( .I1(n15931), .I2(n20628), .O(n19906) );
  MUX2S U25666 ( .A(n20808), .B(n20628), .S(gray_img[65]), .O(n19905) );
  ND2S U25667 ( .I1(n25389), .I2(n20628), .O(n19908) );
  ND2S U25668 ( .I1(n15891), .I2(n20628), .O(n19910) );
  AOI22S U25669 ( .A1(n25103), .A2(n19914), .B1(n25356), .B2(n19913), .O(
        n19915) );
  ND2S U25670 ( .I1(n15937), .I2(n20634), .O(n19917) );
  INV1S U25671 ( .I(gray_img[834]), .O(n22988) );
  ND2S U25672 ( .I1(n15887), .I2(n20634), .O(n19919) );
  INV1S U25673 ( .I(gray_img[835]), .O(n22986) );
  INV1S U25674 ( .I(gray_img[836]), .O(n22984) );
  ND2S U25675 ( .I1(n26828), .I2(n20634), .O(n19923) );
  ND2S U25676 ( .I1(n15888), .I2(n20628), .O(n19925) );
  MUX2S U25677 ( .A(n20808), .B(n20628), .S(gray_img[64]), .O(n19924) );
  ND2S U25678 ( .I1(n15888), .I2(n20634), .O(n19927) );
  INV1S U25679 ( .I(gray_img[832]), .O(n22990) );
  INV1S U25680 ( .I(gray_scale_1[8]), .O(n19928) );
  ND2S U25681 ( .I1(gray_scale_1[9]), .I2(n19928), .O(n19929) );
  ND2S U25682 ( .I1(n19932), .I2(n19929), .O(n30450) );
  INV1S U25683 ( .I(gray_scale_1[7]), .O(n19931) );
  ND2S U25684 ( .I1(n19931), .I2(n19929), .O(n30449) );
  ND2S U25685 ( .I1(n19930), .I2(n30449), .O(n30446) );
  MOAI1S U25686 ( .A1(n19932), .A2(n19931), .B1(n19932), .B2(n19930), .O(
        n30445) );
  INV1S U25687 ( .I(gray_scale_1[6]), .O(n30447) );
  AN2S U25688 ( .I1(n30445), .I2(gray_scale_1[6]), .O(n19933) );
  MOAI1S U25689 ( .A1(n30445), .A2(gray_scale_1[6]), .B1(n30446), .B2(n19933), 
        .O(n19938) );
  ND2S U25690 ( .I1(gray_scale_1[5]), .I2(n19938), .O(n19934) );
  OR2B1S U25691 ( .I1(n19935), .B1(n19934), .O(n30444) );
  OAI12HS U25692 ( .B1(gray_scale_1[5]), .B2(n19935), .A1(n19937), .O(n19941)
         );
  INV1S U25693 ( .I(gray_scale_1[4]), .O(n19940) );
  NR2 U25694 ( .I1(n19940), .I2(n19941), .O(n19939) );
  INV1S U25695 ( .I(n19938), .O(n19936) );
  OAI22S U25696 ( .A1(n19938), .A2(n19937), .B1(n19936), .B2(gray_scale_1[5]), 
        .O(n19944) );
  NR2 U25697 ( .I1(n19939), .I2(n19944), .O(n30443) );
  NR2 U25698 ( .I1(n30443), .I2(n19940), .O(n19942) );
  MOAI1S U25699 ( .A1(n19941), .A2(gray_scale_1[4]), .B1(n19941), .B2(n19942), 
        .O(n19946) );
  INV1S U25700 ( .I(n19942), .O(n19943) );
  ND2S U25701 ( .I1(n19949), .I2(gray_scale_1[3]), .O(n19945) );
  OR2B1S U25702 ( .I1(n19946), .B1(n19945), .O(n30442) );
  OAI12HS U25703 ( .B1(gray_scale_1[3]), .B2(n19946), .A1(n19947), .O(n30439)
         );
  INV1S U25704 ( .I(n19947), .O(n19948) );
  MOAI1S U25705 ( .A1(n19949), .A2(n19948), .B1(n19949), .B2(gray_scale_1[3]), 
        .O(n30438) );
  INV1S U25706 ( .I(gray_scale_1[2]), .O(n30440) );
  AN2S U25707 ( .I1(n30438), .I2(gray_scale_1[2]), .O(n19950) );
  MOAI1S U25708 ( .A1(n30438), .A2(gray_scale_1[2]), .B1(n30439), .B2(n19950), 
        .O(n30436) );
  MOAI1S U25709 ( .A1(n19951), .A2(n30436), .B1(n30436), .B2(gray_scale_1[1]), 
        .O(n19952) );
  ND2S U25710 ( .I1(gray_scale_1_s[0]), .I2(n30452), .O(n19953) );
  ND2S U25711 ( .I1(n19954), .I2(n19953), .O(n13583) );
  ND2S U25712 ( .I1(n15892), .I2(n19955), .O(n19957) );
  ND2S U25713 ( .I1(n15892), .I2(n20449), .O(n19959) );
  ND2S U25714 ( .I1(n20271), .I2(n20550), .O(n19961) );
  ND2S U25715 ( .I1(n20271), .I2(n20463), .O(n19963) );
  ND2S U25716 ( .I1(n25112), .I2(n20528), .O(n19965) );
  ND2S U25717 ( .I1(n15892), .I2(n20504), .O(n19967) );
  ND2S U25718 ( .I1(n20271), .I2(n20596), .O(n19968) );
  ND2S U25719 ( .I1(n25112), .I2(n19970), .O(n19971) );
  ND2S U25720 ( .I1(n25112), .I2(n20608), .O(n19974) );
  ND2S U25721 ( .I1(n19976), .I2(n19975), .O(n14965) );
  MUX2S U25722 ( .A(n20830), .B(n20709), .S(gray_img[1468]), .O(n19977) );
  ND2S U25723 ( .I1(n19980), .I2(n19979), .O(n14980) );
  ND2S U25724 ( .I1(n19982), .I2(n19981), .O(n14964) );
  ND2S U25725 ( .I1(n19984), .I2(n19983), .O(n14990) );
  ND2S U25726 ( .I1(n19986), .I2(n19985), .O(n14974) );
  ND2S U25727 ( .I1(n19988), .I2(n19987), .O(n14950) );
  ND2S U25728 ( .I1(n19990), .I2(n19989), .O(n14966) );
  ND2S U25729 ( .I1(n19992), .I2(n19991), .O(n14998) );
  ND2S U25730 ( .I1(n19994), .I2(n19993), .O(n14982) );
  ND2S U25731 ( .I1(n15890), .I2(n20605), .O(n19995) );
  ND2S U25732 ( .I1(n15890), .I2(n20824), .O(n19997) );
  MUX2S U25733 ( .A(n30005), .B(n20156), .S(gray_img[1830]), .O(n20000) );
  ND2S U25734 ( .I1(n15890), .I2(n20156), .O(n19999) );
  ND2S U25735 ( .I1(n15890), .I2(n20836), .O(n20001) );
  ND2S U25736 ( .I1(n15890), .I2(n20602), .O(n20003) );
  MUX2S U25737 ( .A(n30005), .B(n20202), .S(gray_img[1966]), .O(n20006) );
  ND2S U25738 ( .I1(n15890), .I2(n20202), .O(n20005) );
  ND2S U25739 ( .I1(n15890), .I2(n20827), .O(n20007) );
  ND2S U25740 ( .I1(n15890), .I2(n20814), .O(n20009) );
  MUX2S U25741 ( .A(n30005), .B(n20142), .S(gray_img[1838]), .O(n20012) );
  ND2S U25742 ( .I1(n15890), .I2(n20142), .O(n20011) );
  MUX2S U25743 ( .A(n30005), .B(n20129), .S(gray_img[1310]), .O(n20014) );
  ND2S U25744 ( .I1(n15890), .I2(n20129), .O(n20013) );
  ND2S U25745 ( .I1(n15890), .I2(n20553), .O(n20016) );
  ND2S U25746 ( .I1(n15890), .I2(n20035), .O(n20018) );
  ND2S U25747 ( .I1(n15890), .I2(n20757), .O(n20020) );
  ND2S U25748 ( .I1(n15890), .I2(n20504), .O(n20022) );
  ND2S U25749 ( .I1(n15890), .I2(n20240), .O(n20024) );
  ND2S U25750 ( .I1(n20271), .I2(n20559), .O(n20026) );
  ND2S U25751 ( .I1(n15892), .I2(n20531), .O(n20028) );
  ND2S U25752 ( .I1(n20271), .I2(n20565), .O(n20030) );
  ND2S U25753 ( .I1(n15892), .I2(n20695), .O(n20032) );
  MUX2S U25754 ( .A(n20830), .B(n20695), .S(gray_img[1343]), .O(n20031) );
  ND2S U25755 ( .I1(n15892), .I2(n20547), .O(n20034) );
  ND2S U25756 ( .I1(n25112), .I2(n20035), .O(n20037) );
  ND2S U25757 ( .I1(n15892), .I2(n20731), .O(n20039) );
  ND2S U25758 ( .I1(n15892), .I2(n20427), .O(n20041) );
  MUX2S U25759 ( .A(n20842), .B(n20427), .S(gray_img[1295]), .O(n20040) );
  ND2S U25760 ( .I1(n25112), .I2(n20568), .O(n20043) );
  ND2S U25761 ( .I1(n25112), .I2(n20562), .O(n20045) );
  ND2S U25762 ( .I1(n15892), .I2(n20541), .O(n20047) );
  MUX2S U25763 ( .A(n30005), .B(n20541), .S(gray_img[1783]), .O(n20046) );
  ND2S U25764 ( .I1(n25112), .I2(n20746), .O(n20049) );
  ND2S U25765 ( .I1(n20271), .I2(n20477), .O(n20051) );
  INV1S U25766 ( .I(n25291), .O(n20271) );
  ND2S U25767 ( .I1(n20271), .I2(n20424), .O(n20053) );
  ND2S U25768 ( .I1(n20271), .I2(n20054), .O(n20056) );
  ND2S U25769 ( .I1(n20271), .I2(n20430), .O(n20058) );
  ND2S U25770 ( .I1(n20271), .I2(n20534), .O(n20060) );
  ND2S U25771 ( .I1(n20271), .I2(n20452), .O(n20062) );
  ND2S U25772 ( .I1(n15892), .I2(n20063), .O(n20065) );
  ND2S U25773 ( .I1(n25112), .I2(n20684), .O(n20067) );
  ND2S U25774 ( .I1(n15892), .I2(n20509), .O(n20069) );
  MUX2S U25775 ( .A(n29032), .B(n20509), .S(gray_img[1663]), .O(n20068) );
  ND2S U25776 ( .I1(n20271), .I2(n20725), .O(n20071) );
  MUX2S U25777 ( .A(n20808), .B(n20725), .S(gray_img[1271]), .O(n20070) );
  ND2S U25778 ( .I1(n15892), .I2(n20472), .O(n20073) );
  ND2S U25779 ( .I1(n15892), .I2(n20544), .O(n20075) );
  ND2S U25780 ( .I1(n15892), .I2(n20709), .O(n20077) );
  ND2S U25781 ( .I1(n15892), .I2(n20734), .O(n20079) );
  ND2S U25782 ( .I1(n25112), .I2(n20740), .O(n20081) );
  ND2S U25783 ( .I1(n15892), .I2(n20082), .O(n20084) );
  ND2S U25784 ( .I1(n15892), .I2(n20440), .O(n20086) );
  ND2S U25785 ( .I1(n15892), .I2(n20743), .O(n20088) );
  ND2S U25786 ( .I1(n20271), .I2(n20319), .O(n20090) );
  MUX2S U25787 ( .A(n20808), .B(n20319), .S(gray_img[1807]), .O(n20089) );
  ND2S U25788 ( .I1(n15892), .I2(n20737), .O(n20092) );
  ND2S U25789 ( .I1(n15892), .I2(n20517), .O(n20094) );
  ND2S U25790 ( .I1(n15892), .I2(n20722), .O(n20096) );
  ND2S U25791 ( .I1(n15892), .I2(n20486), .O(n20098) );
  ND2S U25792 ( .I1(n20271), .I2(n20099), .O(n20101) );
  ND2S U25793 ( .I1(n20271), .I2(n20719), .O(n20103) );
  ND2S U25794 ( .I1(n25112), .I2(n20512), .O(n20105) );
  MUX2S U25795 ( .A(n20842), .B(n20512), .S(gray_img[1527]), .O(n20104) );
  ND2S U25796 ( .I1(n15892), .I2(n20525), .O(n20107) );
  MUX2S U25797 ( .A(n30005), .B(n20525), .S(gray_img[1655]), .O(n20106) );
  ND2S U25798 ( .I1(n15892), .I2(n20522), .O(n20109) );
  ND2S U25799 ( .I1(n15892), .I2(n20702), .O(n20111) );
  ND2S U25800 ( .I1(n15892), .I2(n20571), .O(n20113) );
  ND2S U25801 ( .I1(n15892), .I2(n20655), .O(n20115) );
  MUX2S U25802 ( .A(n20808), .B(n20655), .S(gray_img[1279]), .O(n20114) );
  INV1S U25803 ( .I(n25291), .O(n25112) );
  ND2S U25804 ( .I1(n25112), .I2(n20553), .O(n20117) );
  ND2S U25805 ( .I1(n15892), .I2(n20556), .O(n20119) );
  ND2S U25806 ( .I1(n20271), .I2(n20716), .O(n20121) );
  ND2S U25807 ( .I1(n15892), .I2(n20496), .O(n20123) );
  ND2S U25808 ( .I1(n20271), .I2(n20124), .O(n20126) );
  MUX2S U25809 ( .A(n20808), .B(n20124), .S(gray_img[1143]), .O(n20125) );
  ND2S U25810 ( .I1(n25112), .I2(n20728), .O(n20128) );
  MUX2S U25811 ( .A(n30005), .B(n20129), .S(gray_img[1311]), .O(n20131) );
  ND2S U25812 ( .I1(n25112), .I2(n20129), .O(n20130) );
  ND2S U25813 ( .I1(n15892), .I2(n20836), .O(n20132) );
  ND2S U25814 ( .I1(n20271), .I2(n20392), .O(n20134) );
  ND2S U25815 ( .I1(n15892), .I2(n20833), .O(n20136) );
  ND2S U25816 ( .I1(n15892), .I2(n20376), .O(n20138) );
  ND2S U25817 ( .I1(n15892), .I2(n20296), .O(n20140) );
  MUX2S U25818 ( .A(n30005), .B(n20142), .S(gray_img[1839]), .O(n20144) );
  ND2S U25819 ( .I1(n25112), .I2(n20142), .O(n20143) );
  ND2S U25820 ( .I1(n20271), .I2(n20362), .O(n20145) );
  ND2S U25821 ( .I1(n15892), .I2(n20147), .O(n20148) );
  ND2S U25822 ( .I1(n15892), .I2(n20843), .O(n20150) );
  ND2S U25823 ( .I1(n15892), .I2(n20846), .O(n20152) );
  ND2S U25824 ( .I1(n25112), .I2(n20857), .O(n20154) );
  MUX2S U25825 ( .A(n30005), .B(n20156), .S(gray_img[1831]), .O(n20158) );
  ND2S U25826 ( .I1(n25112), .I2(n20156), .O(n20157) );
  ND2S U25827 ( .I1(n25112), .I2(n20159), .O(n20160) );
  ND2S U25828 ( .I1(n15892), .I2(n20379), .O(n20162) );
  ND2S U25829 ( .I1(n15892), .I2(n20787), .O(n20164) );
  ND2S U25830 ( .I1(n15892), .I2(n20591), .O(n20166) );
  ND2S U25831 ( .I1(n25112), .I2(n20293), .O(n20168) );
  ND2S U25832 ( .I1(n15892), .I2(n20839), .O(n20170) );
  ND2S U25833 ( .I1(n15892), .I2(n20583), .O(n20172) );
  ND2S U25834 ( .I1(n20271), .I2(n20862), .O(n20174) );
  ND2S U25835 ( .I1(n15892), .I2(n20811), .O(n20176) );
  ND2S U25836 ( .I1(n15892), .I2(n20814), .O(n20178) );
  ND2S U25837 ( .I1(n15892), .I2(n20821), .O(n20180) );
  ND2S U25838 ( .I1(n20271), .I2(n20365), .O(n20182) );
  ND2S U25839 ( .I1(n20271), .I2(n20184), .O(n20185) );
  ND2S U25840 ( .I1(n15892), .I2(n20827), .O(n20187) );
  MUX2S U25841 ( .A(n30005), .B(n20359), .S(gray_img[1415]), .O(n20190) );
  ND2S U25842 ( .I1(n20271), .I2(n20359), .O(n20189) );
  ND2S U25843 ( .I1(n15892), .I2(n20384), .O(n20191) );
  ND2S U25844 ( .I1(n20271), .I2(n20193), .O(n20194) );
  ND2S U25845 ( .I1(n15892), .I2(n20854), .O(n20196) );
  ND2S U25846 ( .I1(n15892), .I2(n20599), .O(n20198) );
  ND2S U25847 ( .I1(n15892), .I2(n20580), .O(n20200) );
  MUX2S U25848 ( .A(n30005), .B(n20202), .S(gray_img[1967]), .O(n20204) );
  ND2S U25849 ( .I1(n25112), .I2(n20202), .O(n20203) );
  ND2S U25850 ( .I1(n20271), .I2(n20368), .O(n20205) );
  ND2S U25851 ( .I1(n15892), .I2(n20849), .O(n20207) );
  ND2S U25852 ( .I1(n20271), .I2(n20209), .O(n20210) );
  ND2S U25853 ( .I1(n25112), .I2(n20212), .O(n20213) );
  ND2S U25854 ( .I1(n15892), .I2(n20824), .O(n20215) );
  ND2S U25855 ( .I1(n15892), .I2(n20605), .O(n20217) );
  ND2S U25856 ( .I1(n15892), .I2(n20389), .O(n20219) );
  ND2S U25857 ( .I1(n15892), .I2(n20395), .O(n20221) );
  ND2S U25858 ( .I1(n15892), .I2(n20602), .O(n20223) );
  ND2S U25859 ( .I1(n20271), .I2(n20373), .O(n20225) );
  ND2S U25860 ( .I1(n15892), .I2(n25942), .O(n20228) );
  ND2S U25861 ( .I1(n20271), .I2(n20611), .O(n20230) );
  ND2S U25862 ( .I1(n25112), .I2(n20480), .O(n20232) );
  ND2S U25863 ( .I1(n25112), .I2(n20614), .O(n20234) );
  ND2S U25864 ( .I1(n15892), .I2(n20235), .O(n20237) );
  ND2S U25865 ( .I1(n15892), .I2(n20316), .O(n20239) );
  ND2S U25866 ( .I1(n15892), .I2(n20240), .O(n20242) );
  ND2S U25867 ( .I1(n25112), .I2(n20311), .O(n20244) );
  ND2S U25868 ( .I1(n25112), .I2(n20491), .O(n20246) );
  ND2S U25869 ( .I1(n15892), .I2(n20435), .O(n20248) );
  ND2S U25870 ( .I1(n25112), .I2(n20620), .O(n20250) );
  INV1S U25871 ( .I(gray_img[239]), .O(n27406) );
  ND2S U25872 ( .I1(n25112), .I2(n20617), .O(n20252) );
  INV1S U25873 ( .I(gray_img[111]), .O(n25123) );
  ND2S U25874 ( .I1(n15892), .I2(n20623), .O(n20254) );
  ND2S U25875 ( .I1(n15892), .I2(n20255), .O(n20257) );
  ND2S U25876 ( .I1(n25112), .I2(n20483), .O(n20259) );
  MUX2S U25877 ( .A(n30005), .B(n20483), .S(gray_img[455]), .O(n20258) );
  ND2S U25878 ( .I1(n15892), .I2(n20260), .O(n20262) );
  ND2S U25879 ( .I1(n15892), .I2(n20757), .O(n20264) );
  ND2S U25880 ( .I1(n15892), .I2(n20499), .O(n20266) );
  ND2S U25881 ( .I1(n15892), .I2(n20760), .O(n20268) );
  ND2S U25882 ( .I1(n20271), .I2(n20631), .O(n20270) );
  INV1S U25883 ( .I(gray_img[199]), .O(n23614) );
  ND2S U25884 ( .I1(n20271), .I2(n20628), .O(n20273) );
  INV1S U25885 ( .I(gray_img[71]), .O(n23602) );
  ND2S U25886 ( .I1(n25112), .I2(n20274), .O(n20276) );
  MUX2S U25887 ( .A(n30005), .B(n20274), .S(gray_img[623]), .O(n20275) );
  ND2S U25888 ( .I1(n15892), .I2(n20634), .O(n20278) );
  ND2S U25889 ( .I1(n15890), .I2(n20833), .O(n20279) );
  ND2S U25890 ( .I1(n15890), .I2(n20787), .O(n20281) );
  ND2S U25891 ( .I1(n15890), .I2(n20843), .O(n20283) );
  ND2S U25892 ( .I1(n15890), .I2(n20821), .O(n20285) );
  ND2S U25893 ( .I1(n15890), .I2(n20857), .O(n20287) );
  ND2S U25894 ( .I1(n15890), .I2(n20811), .O(n20289) );
  ND2S U25895 ( .I1(n15890), .I2(n20854), .O(n20291) );
  ND2S U25896 ( .I1(n15890), .I2(n20293), .O(n20294) );
  ND2S U25897 ( .I1(n15890), .I2(n20296), .O(n20297) );
  ND2S U25898 ( .I1(n15890), .I2(n20583), .O(n20299) );
  ND2S U25899 ( .I1(n15890), .I2(n20760), .O(n20302) );
  ND2S U25900 ( .I1(n15890), .I2(n20695), .O(n20304) );
  MUX2S U25901 ( .A(n20830), .B(n20695), .S(gray_img[1342]), .O(n20303) );
  ND2S U25902 ( .I1(n15890), .I2(n20709), .O(n20306) );
  MUX2S U25903 ( .A(n20830), .B(n20709), .S(gray_img[1470]), .O(n20305) );
  ND2S U25904 ( .I1(n15890), .I2(n20655), .O(n20308) );
  MUX2S U25905 ( .A(n20808), .B(n20655), .S(gray_img[1278]), .O(n20307) );
  ND2S U25906 ( .I1(n15890), .I2(n20559), .O(n20310) );
  ND2S U25907 ( .I1(n15890), .I2(n20311), .O(n20313) );
  ND2S U25908 ( .I1(n15890), .I2(n20531), .O(n20315) );
  ND2S U25909 ( .I1(n15890), .I2(n20316), .O(n20318) );
  ND2S U25910 ( .I1(n15890), .I2(n20319), .O(n20321) );
  MOAI1S U25911 ( .A1(n20322), .A2(n25062), .B1(n25193), .B2(n25061), .O(
        n20323) );
  MUX2S U25912 ( .A(n30005), .B(n20586), .S(gray_img[1957]), .O(n20325) );
  ND2S U25913 ( .I1(n26828), .I2(n20586), .O(n20324) );
  ND2S U25914 ( .I1(n20325), .I2(n20324), .O(n15088) );
  MUX2S U25915 ( .A(n30005), .B(n20586), .S(gray_img[1956]), .O(n20327) );
  MUX2S U25916 ( .A(n30005), .B(n20586), .S(gray_img[1959]), .O(n20329) );
  ND2S U25917 ( .I1(n25112), .I2(n20586), .O(n20328) );
  MUX2S U25918 ( .A(n30005), .B(n20586), .S(gray_img[1955]), .O(n20331) );
  ND2S U25919 ( .I1(n15887), .I2(n20586), .O(n20330) );
  ND2S U25920 ( .I1(n20331), .I2(n20330), .O(n14689) );
  MUX2S U25921 ( .A(n30005), .B(n20586), .S(gray_img[1954]), .O(n20333) );
  ND2S U25922 ( .I1(n15883), .I2(n20586), .O(n20332) );
  ND2S U25923 ( .I1(n20333), .I2(n20332), .O(n14489) );
  MOAI1S U25924 ( .A1(n20334), .A2(n25066), .B1(n25272), .B2(n25065), .O(
        n20335) );
  ND2S U25925 ( .I1(n15891), .I2(n20354), .O(n20336) );
  ND2S U25926 ( .I1(n20337), .I2(n20336), .O(n15106) );
  ND2S U25927 ( .I1(n15892), .I2(n20354), .O(n20340) );
  ND2S U25928 ( .I1(n15883), .I2(n20354), .O(n20342) );
  ND2S U25929 ( .I1(n20343), .I2(n20342), .O(n14507) );
  ND2S U25930 ( .I1(n15887), .I2(n20354), .O(n20344) );
  ND2S U25931 ( .I1(n20345), .I2(n20344), .O(n14707) );
  MUX2S U25932 ( .A(n30005), .B(n20586), .S(gray_img[1958]), .O(n20347) );
  ND2S U25933 ( .I1(n15890), .I2(n20586), .O(n20346) );
  MUX2S U25934 ( .A(n30005), .B(n20586), .S(gray_img[1952]), .O(n20349) );
  ND2S U25935 ( .I1(n15888), .I2(n20586), .O(n20348) );
  ND2S U25936 ( .I1(n20349), .I2(n20348), .O(n13832) );
  ND2S U25937 ( .I1(n15890), .I2(n20354), .O(n20350) );
  ND2S U25938 ( .I1(n15888), .I2(n20354), .O(n20352) );
  ND2S U25939 ( .I1(n20353), .I2(n20352), .O(n13857) );
  ND2S U25940 ( .I1(n20356), .I2(n20355), .O(n14306) );
  ND2S U25941 ( .I1(n25389), .I2(n20849), .O(n20357) );
  ND2S U25942 ( .I1(n25444), .I2(n20359), .O(n20360) );
  ND2S U25943 ( .I1(n25448), .I2(n20362), .O(n20363) );
  ND2S U25944 ( .I1(n25389), .I2(n20365), .O(n20366) );
  ND2S U25945 ( .I1(n15890), .I2(n20368), .O(n20369) );
  ND2S U25946 ( .I1(n20370), .I2(n20369), .O(n15396) );
  ND2S U25947 ( .I1(n25444), .I2(n20862), .O(n20371) );
  ND2S U25948 ( .I1(n25448), .I2(n20373), .O(n20374) );
  ND2S U25949 ( .I1(n25444), .I2(n20376), .O(n20377) );
  ND2S U25950 ( .I1(n20378), .I2(n20377), .O(n15304) );
  ND2S U25951 ( .I1(n25389), .I2(n20379), .O(n20380) );
  ND2S U25952 ( .I1(n20381), .I2(n20380), .O(n15380) );
  ND2S U25953 ( .I1(n25448), .I2(n20599), .O(n20382) );
  ND2S U25954 ( .I1(n15890), .I2(n20384), .O(n20385) );
  ND2S U25955 ( .I1(n20386), .I2(n20385), .O(n15403) );
  ND2S U25956 ( .I1(n25389), .I2(n20839), .O(n20387) );
  ND2S U25957 ( .I1(n25444), .I2(n20389), .O(n20390) );
  ND2S U25958 ( .I1(n25389), .I2(n20392), .O(n20393) );
  ND2S U25959 ( .I1(n25444), .I2(n20395), .O(n20396) );
  ND2S U25960 ( .I1(n25448), .I2(n20591), .O(n20398) );
  ND2S U25961 ( .I1(n20399), .I2(n20398), .O(n15432) );
  ND2S U25962 ( .I1(n25448), .I2(n20846), .O(n20400) );
  ND2S U25963 ( .I1(n15890), .I2(n20544), .O(n20403) );
  ND2S U25964 ( .I1(n15890), .I2(n20737), .O(n20405) );
  ND2S U25965 ( .I1(n15890), .I2(n20556), .O(n20407) );
  ND2S U25966 ( .I1(n15890), .I2(n20740), .O(n20409) );
  ND2S U25967 ( .I1(n15890), .I2(n20731), .O(n20411) );
  ND2S U25968 ( .I1(n25448), .I2(n25942), .O(n20413) );
  MUX2S U25969 ( .A(n30005), .B(n25942), .S(gray_img[2038]), .O(n20412) );
  ND2S U25970 ( .I1(n20413), .I2(n20412), .O(n15274) );
  ND2S U25971 ( .I1(n25444), .I2(n20684), .O(n20415) );
  ND2S U25972 ( .I1(n15890), .I2(n20608), .O(n20417) );
  ND2S U25973 ( .I1(n15890), .I2(n20746), .O(n20419) );
  ND2S U25974 ( .I1(n25448), .I2(n20517), .O(n20421) );
  ND2S U25975 ( .I1(n20421), .I2(n20420), .O(n15354) );
  ND2S U25976 ( .I1(n25444), .I2(n20614), .O(n20423) );
  MUX2S U25977 ( .A(n30005), .B(n20614), .S(gray_img[2046]), .O(n20422) );
  ND2S U25978 ( .I1(n20423), .I2(n20422), .O(n15273) );
  ND2S U25979 ( .I1(n15890), .I2(n20424), .O(n20426) );
  ND2S U25980 ( .I1(n25448), .I2(n20427), .O(n20429) );
  ND2S U25981 ( .I1(n15890), .I2(n20430), .O(n20432) );
  ND2S U25982 ( .I1(n25444), .I2(n20702), .O(n20434) );
  ND2S U25983 ( .I1(n20434), .I2(n20433), .O(n15376) );
  ND2S U25984 ( .I1(n25448), .I2(n20435), .O(n20437) );
  ND2S U25985 ( .I1(n15890), .I2(n20547), .O(n20439) );
  ND2S U25986 ( .I1(n25444), .I2(n20440), .O(n20442) );
  ND2S U25987 ( .I1(n20442), .I2(n20441), .O(n15339) );
  ND2S U25988 ( .I1(n25389), .I2(n20743), .O(n20444) );
  ND2S U25989 ( .I1(n20444), .I2(n20443), .O(n15392) );
  ND2S U25990 ( .I1(n25448), .I2(n20611), .O(n20446) );
  ND2S U25991 ( .I1(n15890), .I2(n20541), .O(n20448) );
  ND2S U25992 ( .I1(n15890), .I2(n20449), .O(n20451) );
  ND2S U25993 ( .I1(n25389), .I2(n20452), .O(n20454) );
  ND2S U25994 ( .I1(n25444), .I2(n20722), .O(n20456) );
  ND2S U25995 ( .I1(n15890), .I2(n20634), .O(n20458) );
  INV1S U25996 ( .I(gray_img[838]), .O(n22971) );
  ND2S U25997 ( .I1(n25444), .I2(n20568), .O(n20460) );
  ND2S U25998 ( .I1(n25448), .I2(n20509), .O(n20462) );
  MUX2S U25999 ( .A(n29032), .B(n20509), .S(gray_img[1662]), .O(n20461) );
  ND2S U26000 ( .I1(n25389), .I2(n20463), .O(n20465) );
  MUX2S U26001 ( .A(n29032), .B(n20463), .S(gray_img[1646]), .O(n20464) );
  ND2S U26002 ( .I1(n20465), .I2(n20464), .O(n15323) );
  ND2S U26003 ( .I1(n25389), .I2(n20565), .O(n20467) );
  ND2S U26004 ( .I1(n25444), .I2(n20534), .O(n20469) );
  ND2S U26005 ( .I1(n25448), .I2(n20716), .O(n20471) );
  ND2S U26006 ( .I1(n20471), .I2(n20470), .O(n15385) );
  ND2S U26007 ( .I1(n15890), .I2(n20472), .O(n20474) );
  ND2S U26008 ( .I1(n20474), .I2(n20473), .O(n15433) );
  ND2S U26009 ( .I1(n25448), .I2(n20512), .O(n20476) );
  MUX2S U26010 ( .A(n20830), .B(n20512), .S(gray_img[1526]), .O(n20475) );
  ND2S U26011 ( .I1(n25389), .I2(n20477), .O(n20479) );
  ND2S U26012 ( .I1(n25444), .I2(n20480), .O(n20482) );
  ND2S U26013 ( .I1(n25444), .I2(n20483), .O(n20485) );
  ND2S U26014 ( .I1(n25448), .I2(n20486), .O(n20488) );
  ND2S U26015 ( .I1(n25389), .I2(n20522), .O(n20490) );
  ND2S U26016 ( .I1(n20490), .I2(n20489), .O(n15442) );
  ND2S U26017 ( .I1(n25448), .I2(n20491), .O(n20493) );
  ND2S U26018 ( .I1(n15890), .I2(n20620), .O(n20495) );
  INV1S U26019 ( .I(gray_img[238]), .O(n27405) );
  ND2S U26020 ( .I1(n20495), .I2(n20494), .O(n15451) );
  ND2S U26021 ( .I1(n25444), .I2(n20496), .O(n20498) );
  ND2S U26022 ( .I1(n20498), .I2(n20497), .O(n15449) );
  ND2S U26023 ( .I1(n25389), .I2(n20499), .O(n20501) );
  ND2S U26024 ( .I1(n25448), .I2(n20617), .O(n20503) );
  INV1S U26025 ( .I(gray_img[110]), .O(n27401) );
  ND2S U26026 ( .I1(n20506), .I2(n20505), .O(n14300) );
  ND2S U26027 ( .I1(n20508), .I2(n20507), .O(n14724) );
  ND2S U26028 ( .I1(n20511), .I2(n20510), .O(n14526) );
  ND2S U26029 ( .I1(n20514), .I2(n20513), .O(n14743) );
  ND2S U26030 ( .I1(n20516), .I2(n20515), .O(n14831) );
  ND2S U26031 ( .I1(n20519), .I2(n20518), .O(n14759) );
  ND2S U26032 ( .I1(n20521), .I2(n20520), .O(n14540) );
  ND2S U26033 ( .I1(n20524), .I2(n20523), .O(n14847) );
  ND2S U26034 ( .I1(n20527), .I2(n20526), .O(n14527) );
  MUX2S U26035 ( .A(n29032), .B(n20528), .S(gray_img[1601]), .O(n20529) );
  ND2S U26036 ( .I1(n20530), .I2(n20529), .O(n14332) );
  ND2S U26037 ( .I1(n20533), .I2(n20532), .O(n14524) );
  ND2S U26038 ( .I1(n20536), .I2(n20535), .O(n14631) );
  ND2S U26039 ( .I1(n20538), .I2(n20537), .O(n14815) );
  ND2S U26040 ( .I1(n20540), .I2(n20539), .O(n14807) );
  ND2S U26041 ( .I1(n20543), .I2(n20542), .O(n14511) );
  ND2S U26042 ( .I1(n20546), .I2(n20545), .O(n14295) );
  ND2S U26043 ( .I1(n20549), .I2(n20548), .O(n14510) );
  ND2S U26044 ( .I1(n20552), .I2(n20551), .O(n14740) );
  ND2S U26045 ( .I1(n20555), .I2(n20554), .O(n14788) );
  ND2S U26046 ( .I1(n20558), .I2(n20557), .O(n14742) );
  ND2S U26047 ( .I1(n20561), .I2(n20560), .O(n14615) );
  ND2S U26048 ( .I1(n20564), .I2(n20563), .O(n14607) );
  ND2S U26049 ( .I1(n20567), .I2(n20566), .O(n14429) );
  ND2S U26050 ( .I1(n20570), .I2(n20569), .O(n14421) );
  ND2S U26051 ( .I1(n20573), .I2(n20572), .O(n14758) );
  ND2S U26052 ( .I1(n20575), .I2(n20574), .O(n14538) );
  ND2S U26053 ( .I1(n20577), .I2(n20576), .O(n14725) );
  ND2S U26054 ( .I1(n20579), .I2(n20578), .O(n14523) );
  ND2S U26055 ( .I1(n20582), .I2(n20581), .O(n14412) );
  ND2S U26056 ( .I1(n20585), .I2(n20584), .O(n14525) );
  MUX2S U26057 ( .A(n30005), .B(n20586), .S(gray_img[1953]), .O(n20588) );
  ND2S U26058 ( .I1(n20588), .I2(n20587), .O(n14288) );
  MUX2S U26059 ( .A(n29032), .B(n20599), .S(gray_img[1690]), .O(n20590) );
  ND2S U26060 ( .I1(n20590), .I2(n20589), .O(n14522) );
  ND2S U26061 ( .I1(n20593), .I2(n20592), .O(n14436) );
  ND2S U26062 ( .I1(n20595), .I2(n20594), .O(n14739) );
  ND2S U26063 ( .I1(n20598), .I2(n20597), .O(n14738) );
  ND2S U26064 ( .I1(n20601), .I2(n20600), .O(n14722) );
  ND2S U26065 ( .I1(n20604), .I2(n20603), .O(n14539) );
  ND2S U26066 ( .I1(n20607), .I2(n20606), .O(n14723) );
  MUX2S U26067 ( .A(n30005), .B(n20608), .S(gray_img[2025]), .O(n20609) );
  ND2S U26068 ( .I1(n20610), .I2(n20609), .O(n14279) );
  ND2S U26069 ( .I1(n20613), .I2(n20612), .O(n14600) );
  MUX2S U26070 ( .A(n30005), .B(n20614), .S(gray_img[2041]), .O(n20615) );
  ND2S U26071 ( .I1(n20616), .I2(n20615), .O(n14277) );
  ND2S U26072 ( .I1(n20619), .I2(n20618), .O(n14463) );
  ND2S U26073 ( .I1(n20622), .I2(n20621), .O(n14455) );
  MUX2S U26074 ( .A(n20808), .B(n20628), .S(gray_img[66]), .O(n20626) );
  MUX2S U26075 ( .A(n20808), .B(n20628), .S(gray_img[67]), .O(n20629) );
  MUX2S U26076 ( .A(n20634), .B(n20830), .S(intadd_99_CI), .O(n20635) );
  ND2S U26077 ( .I1(n20638), .I2(n20637), .O(n14317) );
  ND2S U26078 ( .I1(n20640), .I2(n20639), .O(n14781) );
  ND2S U26079 ( .I1(n20642), .I2(n20641), .O(n14348) );
  ND2S U26080 ( .I1(n20644), .I2(n20643), .O(n14565) );
  ND2S U26081 ( .I1(n20646), .I2(n20645), .O(n14790) );
  ND2S U26082 ( .I1(n20648), .I2(n20647), .O(n14774) );
  ND2S U26083 ( .I1(n20650), .I2(n20649), .O(n14549) );
  ND2S U26084 ( .I1(n20652), .I2(n20651), .O(n14776) );
  ND2S U26085 ( .I1(n20654), .I2(n20653), .O(n14574) );
  ND2S U26086 ( .I1(n20657), .I2(n20656), .O(n14373) );
  ND2S U26087 ( .I1(n20659), .I2(n20658), .O(n14560) );
  ND2S U26088 ( .I1(n20661), .I2(n20660), .O(n14575) );
  ND2S U26089 ( .I1(n20663), .I2(n20662), .O(n14576) );
  ND2S U26090 ( .I1(n20665), .I2(n20664), .O(n14534) );
  ND2S U26091 ( .I1(n20667), .I2(n20666), .O(n14792) );
  ND2S U26092 ( .I1(n20669), .I2(n20668), .O(n14797) );
  ND2S U26093 ( .I1(n20671), .I2(n20670), .O(n14502) );
  ND2S U26094 ( .I1(n20673), .I2(n20672), .O(n14285) );
  MUX2S U26095 ( .A(n20830), .B(n20709), .S(gray_img[1467]), .O(n20674) );
  ND2S U26096 ( .I1(n20675), .I2(n20674), .O(n14750) );
  ND2S U26097 ( .I1(n20677), .I2(n20676), .O(n14349) );
  ND2S U26098 ( .I1(n20679), .I2(n20678), .O(n14389) );
  ND2S U26099 ( .I1(n20681), .I2(n20680), .O(n14365) );
  ND2S U26100 ( .I1(n20683), .I2(n20682), .O(n14566) );
  ND2S U26101 ( .I1(n20686), .I2(n20685), .O(n14749) );
  ND2S U26102 ( .I1(n20688), .I2(n20687), .O(n14391) );
  ND2S U26103 ( .I1(n20690), .I2(n20689), .O(n14333) );
  ND2S U26104 ( .I1(n20692), .I2(n20691), .O(n14775) );
  ND2S U26105 ( .I1(n20694), .I2(n20693), .O(n14581) );
  ND2S U26106 ( .I1(n20697), .I2(n20696), .O(n14766) );
  ND2S U26107 ( .I1(n20699), .I2(n20698), .O(n14765) );
  ND2S U26108 ( .I1(n20701), .I2(n20700), .O(n14301) );
  ND2S U26109 ( .I1(n20704), .I2(n20703), .O(n14380) );
  ND2S U26110 ( .I1(n20706), .I2(n20705), .O(n14760) );
  ND2S U26111 ( .I1(n20708), .I2(n20707), .O(n14396) );
  MUX2S U26112 ( .A(n20830), .B(n20709), .S(gray_img[1466]), .O(n20710) );
  ND2S U26113 ( .I1(n20711), .I2(n20710), .O(n14550) );
  ND2S U26114 ( .I1(n20713), .I2(n20712), .O(n14718) );
  ND2S U26115 ( .I1(n20715), .I2(n20714), .O(n14486) );
  ND2S U26116 ( .I1(n20718), .I2(n20717), .O(n14590) );
  ND2S U26117 ( .I1(n20721), .I2(n20720), .O(n14375) );
  ND2S U26118 ( .I1(n20724), .I2(n20723), .O(n14359) );
  ND2S U26119 ( .I1(n20727), .I2(n20726), .O(n14374) );
  MUX2S U26120 ( .A(n20830), .B(n20728), .S(gray_img[1130]), .O(n20729) );
  ND2S U26121 ( .I1(n20730), .I2(n20729), .O(n14592) );
  ND2S U26122 ( .I1(n20733), .I2(n20732), .O(n14734) );
  ND2S U26123 ( .I1(n20736), .I2(n20735), .O(n14364) );
  ND2S U26124 ( .I1(n20739), .I2(n20738), .O(n14518) );
  ND2S U26125 ( .I1(n20742), .I2(n20741), .O(n14702) );
  ND2S U26126 ( .I1(n20745), .I2(n20744), .O(n14597) );
  ND2S U26127 ( .I1(n20748), .I2(n20747), .O(n14686) );
  ND2S U26128 ( .I1(n20764), .I2(n20763), .O(n14302) );
  ND2S U26129 ( .I1(n20766), .I2(n20765), .O(n14286) );
  ND2S U26130 ( .I1(n20768), .I2(n20767), .O(n14318) );
  ND2S U26131 ( .I1(n20770), .I2(n20769), .O(n14319) );
  ND2S U26132 ( .I1(n20772), .I2(n20771), .O(n14334) );
  ND2S U26133 ( .I1(n20774), .I2(n20773), .O(n14551) );
  ND2S U26134 ( .I1(n20776), .I2(n20775), .O(n14351) );
  ND2S U26135 ( .I1(n20778), .I2(n20777), .O(n14552) );
  MUX2S U26136 ( .A(n30050), .B(n20811), .S(gray_img[1442]), .O(n20780) );
  ND2S U26137 ( .I1(n20780), .I2(n20779), .O(n14553) );
  ND2S U26138 ( .I1(n20782), .I2(n20781), .O(n14799) );
  ND2S U26139 ( .I1(n20784), .I2(n20783), .O(n14567) );
  ND2S U26140 ( .I1(n20786), .I2(n20785), .O(n14783) );
  ND2S U26141 ( .I1(n20789), .I2(n20788), .O(n14320) );
  ND2S U26142 ( .I1(n20791), .I2(n20790), .O(n14568) );
  ND2S U26143 ( .I1(n20793), .I2(n20792), .O(n14487) );
  ND2S U26144 ( .I1(n20795), .I2(n20794), .O(n14720) );
  ND2S U26145 ( .I1(n20797), .I2(n20796), .O(n14537) );
  ND2S U26146 ( .I1(n20799), .I2(n20798), .O(n14569) );
  ND2S U26147 ( .I1(n20801), .I2(n20800), .O(n14769) );
  ND2S U26148 ( .I1(n20803), .I2(n20802), .O(n14535) );
  ND2S U26149 ( .I1(n20805), .I2(n20804), .O(n14768) );
  ND2S U26150 ( .I1(n20807), .I2(n20806), .O(n14767) );
  ND2S U26151 ( .I1(n20810), .I2(n20809), .O(n14352) );
  MUX2S U26152 ( .A(n30005), .B(n20811), .S(gray_img[1443]), .O(n20813) );
  ND2S U26153 ( .I1(n20813), .I2(n20812), .O(n14753) );
  ND2S U26154 ( .I1(n20816), .I2(n20815), .O(n14752) );
  ND2S U26155 ( .I1(n20818), .I2(n20817), .O(n14751) );
  ND2S U26156 ( .I1(n20820), .I2(n20819), .O(n14583) );
  ND2S U26157 ( .I1(n20823), .I2(n20822), .O(n14350) );
  ND2S U26158 ( .I1(n20826), .I2(n20825), .O(n14737) );
  ND2S U26159 ( .I1(n20829), .I2(n20828), .O(n14520) );
  ND2S U26160 ( .I1(n20832), .I2(n20831), .O(n14519) );
  ND2S U26161 ( .I1(n20835), .I2(n20834), .O(n14366) );
  ND2S U26162 ( .I1(n20838), .I2(n20837), .O(n14367) );
  ND2S U26163 ( .I1(n20841), .I2(n20840), .O(n14735) );
  ND2S U26164 ( .I1(n20845), .I2(n20844), .O(n14368) );
  ND2S U26165 ( .I1(n20848), .I2(n20847), .O(n14719) );
  ND2S U26166 ( .I1(n20851), .I2(n20850), .O(n14687) );
  ND2S U26167 ( .I1(n20853), .I2(n20852), .O(n14398) );
  ND2S U26168 ( .I1(n20856), .I2(n20855), .O(n14599) );
  ND2S U26169 ( .I1(n20859), .I2(n20858), .O(n14382) );
  ND2S U26170 ( .I1(n20861), .I2(n20860), .O(n14703) );
  ND2S U26171 ( .I1(n20864), .I2(n20863), .O(n14503) );
  MOAI1S U26172 ( .A1(n20865), .A2(n25054), .B1(n25216), .B2(n25053), .O(
        n20866) );
  ND2S U26173 ( .I1(n20868), .I2(n20867), .O(n14741) );
  ND2S U26174 ( .I1(n20870), .I2(n20869), .O(n14541) );
  ND2S U26175 ( .I1(n15891), .I2(n20881), .O(n20871) );
  ND2S U26176 ( .I1(n20872), .I2(n20871), .O(n15140) );
  ND2S U26177 ( .I1(n15892), .I2(n20881), .O(n20875) );
  ND2S U26178 ( .I1(n15884), .I2(n20881), .O(n20877) );
  ND2S U26179 ( .I1(n20878), .I2(n20877), .O(n14340) );
  ND2S U26180 ( .I1(n15890), .I2(n20881), .O(n20879) );
  ND2S U26181 ( .I1(n15888), .I2(n20881), .O(n20882) );
  ND2S U26182 ( .I1(n20883), .I2(n20882), .O(n13923) );
  AOI22S U26183 ( .A1(n25372), .A2(n25086), .B1(n25370), .B2(n25085), .O(
        n20884) );
  OA12S U26184 ( .B1(gray_img[415]), .B2(n29427), .A1(n28728), .O(n20885) );
  MOAI1S U26185 ( .A1(n28728), .A2(gray_img[415]), .B1(n25291), .B2(n20885), 
        .O(n20888) );
  INV1S U26186 ( .I(gray_img[831]), .O(n25080) );
  INV1S U26187 ( .I(gray_img[959]), .O(n26123) );
  ND2S U26188 ( .I1(n25080), .I2(n26123), .O(n26132) );
  INV1S U26189 ( .I(n26132), .O(n20886) );
  NR2 U26190 ( .I1(gray_img[823]), .I2(gray_img[951]), .O(n26131) );
  AO12S U26191 ( .B1(n20886), .B2(n26131), .A1(n29680), .O(n20887) );
  ND2S U26192 ( .I1(n20888), .I2(n20887), .O(n15467) );
  AOI22S U26193 ( .A1(n25195), .A2(n25274), .B1(n25333), .B2(n25272), .O(
        n20889) );
  OA12S U26194 ( .B1(gray_img[535]), .B2(n29427), .A1(n29044), .O(n20890) );
  MOAI1S U26195 ( .A1(n29044), .A2(gray_img[535]), .B1(n25291), .B2(n20890), 
        .O(n20894) );
  INV1S U26196 ( .I(gray_img[1071]), .O(n20891) );
  INV1S U26197 ( .I(gray_img[1199]), .O(n23032) );
  ND2S U26198 ( .I1(n20891), .I2(n23032), .O(n23041) );
  INV1S U26199 ( .I(n23041), .O(n20892) );
  NR2 U26200 ( .I1(gray_img[1191]), .I2(gray_img[1063]), .O(n23040) );
  AO12S U26201 ( .B1(n20892), .B2(n23040), .A1(n29680), .O(n20893) );
  ND2S U26202 ( .I1(n20894), .I2(n20893), .O(n14048) );
  AOI22S U26203 ( .A1(n25103), .A2(n25245), .B1(n25356), .B2(n25244), .O(
        n20895) );
  OA12S U26204 ( .B1(gray_img[815]), .B2(n29427), .A1(n25605), .O(n20896) );
  MOAI1S U26205 ( .A1(n25605), .A2(gray_img[815]), .B1(n25291), .B2(n20896), 
        .O(n20900) );
  INV1S U26206 ( .I(gray_img[1759]), .O(n20897) );
  INV1S U26207 ( .I(gray_img[1631]), .O(n25537) );
  ND2S U26208 ( .I1(n20897), .I2(n25537), .O(n25546) );
  INV1S U26209 ( .I(n25546), .O(n20898) );
  NR2 U26210 ( .I1(gray_img[1623]), .I2(gray_img[1751]), .O(n25545) );
  AO12S U26211 ( .B1(n20898), .B2(n25545), .A1(n29680), .O(n20899) );
  ND2S U26212 ( .I1(n20900), .I2(n20899), .O(n13872) );
  AOI22S U26213 ( .A1(n25162), .A2(n25245), .B1(n25361), .B2(n25244), .O(
        n20901) );
  OA12S U26214 ( .B1(gray_img[303]), .B2(n29427), .A1(n27114), .O(n20902) );
  MOAI1S U26215 ( .A1(n27114), .A2(gray_img[303]), .B1(n25291), .B2(n20902), 
        .O(n20906) );
  INV1S U26216 ( .I(gray_img[727]), .O(n20903) );
  ND2S U26217 ( .I1(n20903), .I2(n27025), .O(n27046) );
  INV1S U26218 ( .I(n27046), .O(n20904) );
  NR2 U26219 ( .I1(gray_img[607]), .I2(gray_img[735]), .O(n27045) );
  AO12S U26220 ( .B1(n20904), .B2(n27045), .A1(n29680), .O(n20905) );
  ND2S U26221 ( .I1(n20906), .I2(n20905), .O(n14153) );
  AOI22S U26222 ( .A1(n25218), .A2(n25372), .B1(n25216), .B2(n25370), .O(
        n20907) );
  OA12S U26223 ( .B1(gray_img[391]), .B2(n29427), .A1(n30103), .O(n20908) );
  MOAI1S U26224 ( .A1(n30103), .A2(gray_img[391]), .B1(n25291), .B2(n20908), 
        .O(n20911) );
  INV1S U26225 ( .I(gray_img[783]), .O(n25094) );
  ND2S U26226 ( .I1(n25094), .I2(n29616), .O(n29637) );
  INV1S U26227 ( .I(n29637), .O(n20909) );
  NR2 U26228 ( .I1(gray_img[903]), .I2(gray_img[775]), .O(n29636) );
  AO12S U26229 ( .B1(n20909), .B2(n29636), .A1(n29680), .O(n20910) );
  ND2S U26230 ( .I1(n20911), .I2(n20910), .O(n13631) );
  AOI22S U26231 ( .A1(n25326), .A2(n25217), .B1(n25325), .B2(n25347), .O(
        n20912) );
  OA12S U26232 ( .B1(gray_img[911]), .B2(n29427), .A1(n29598), .O(n20913) );
  MOAI1S U26233 ( .A1(n29598), .A2(gray_img[911]), .B1(n25291), .B2(n20913), 
        .O(n20917) );
  INV1S U26234 ( .I(gray_img[1823]), .O(n20914) );
  INV1S U26235 ( .I(gray_img[1951]), .O(n29516) );
  ND2S U26236 ( .I1(n20914), .I2(n29516), .O(n29523) );
  INV1S U26237 ( .I(n29523), .O(n20915) );
  NR2 U26238 ( .I1(gray_img[1943]), .I2(gray_img[1815]), .O(n29522) );
  AO12S U26239 ( .B1(n20915), .B2(n29522), .A1(n29680), .O(n20916) );
  ND2S U26240 ( .I1(n20917), .I2(n20916), .O(n13833) );
  AOI22S U26241 ( .A1(n25246), .A2(n25326), .B1(n25257), .B2(n25325), .O(
        n20918) );
  OA12S U26242 ( .B1(gray_img[143]), .B2(n29427), .A1(n28840), .O(n20919) );
  MOAI1S U26243 ( .A1(n28840), .A2(gray_img[143]), .B1(n25291), .B2(n20919), 
        .O(n20923) );
  INV1S U26244 ( .I(gray_img[279]), .O(n20920) );
  ND2S U26245 ( .I1(n20920), .I2(n28746), .O(n28773) );
  INV1S U26246 ( .I(n28773), .O(n20921) );
  NR2 U26247 ( .I1(gray_img[415]), .I2(gray_img[287]), .O(n28772) );
  AO12S U26248 ( .B1(n20921), .B2(n28772), .A1(n29680), .O(n20922) );
  ND2S U26249 ( .I1(n20923), .I2(n20922), .O(n15466) );
  AOI22S U26250 ( .A1(n25195), .A2(n25283), .B1(n25333), .B2(n25282), .O(
        n20924) );
  OA12S U26251 ( .B1(gray_img[575]), .B2(n29427), .A1(n23493), .O(n20925) );
  MOAI1S U26252 ( .A1(gray_img[575]), .A2(n23493), .B1(n25291), .B2(n20925), 
        .O(n20929) );
  INV1S U26253 ( .I(gray_img[1151]), .O(n20926) );
  INV1S U26254 ( .I(gray_img[1279]), .O(n23323) );
  ND2S U26255 ( .I1(n20926), .I2(n23323), .O(n23332) );
  INV1S U26256 ( .I(n23332), .O(n20927) );
  NR2 U26257 ( .I1(gray_img[1143]), .I2(gray_img[1271]), .O(n23331) );
  AO12S U26258 ( .B1(n20927), .B2(n23331), .A1(n29680), .O(n20928) );
  ND2S U26259 ( .I1(n20929), .I2(n20928), .O(n14003) );
  AOI22S U26260 ( .A1(n25373), .A2(n25162), .B1(n25371), .B2(n25361), .O(
        n20930) );
  OA12S U26261 ( .B1(gray_img[311]), .B2(n29427), .A1(n26322), .O(n20931) );
  MOAI1S U26262 ( .A1(n26322), .A2(gray_img[311]), .B1(n25291), .B2(n20931), 
        .O(n20934) );
  OR2S U26263 ( .I1(gray_img[615]), .I2(gray_img[743]), .O(n26202) );
  INV1S U26264 ( .I(n26202), .O(n20932) );
  NR2 U26265 ( .I1(gray_img[623]), .I2(gray_img[751]), .O(n26203) );
  AO12S U26266 ( .B1(n20932), .B2(n26203), .A1(n29680), .O(n20933) );
  ND2S U26267 ( .I1(n20934), .I2(n20933), .O(n14144) );
  AOI22S U26268 ( .A1(n25162), .A2(n25274), .B1(n25361), .B2(n25272), .O(
        n20935) );
  OA12S U26269 ( .B1(gray_img[279]), .B2(n29427), .A1(n28707), .O(n20936) );
  MOAI1S U26270 ( .A1(n28707), .A2(gray_img[279]), .B1(n25291), .B2(n20936), 
        .O(n20939) );
  INV1S U26271 ( .I(gray_img[679]), .O(n25210) );
  ND2S U26272 ( .I1(n25210), .I2(n28632), .O(n28641) );
  INV1S U26273 ( .I(n28641), .O(n20937) );
  NR2 U26274 ( .I1(gray_img[559]), .I2(gray_img[687]), .O(n28640) );
  AO12S U26275 ( .B1(n20937), .B2(n28640), .A1(n29680), .O(n20938) );
  ND2S U26276 ( .I1(n20939), .I2(n20938), .O(n13674) );
  AOI22S U26277 ( .A1(n25086), .A2(n25217), .B1(n25085), .B2(n25347), .O(
        n20940) );
  OA12S U26278 ( .B1(gray_img[927]), .B2(n29427), .A1(n23195), .O(n20941) );
  MOAI1S U26279 ( .A1(n23195), .A2(gray_img[927]), .B1(n25291), .B2(n20941), 
        .O(n20945) );
  INV1S U26280 ( .I(gray_img[1847]), .O(n20942) );
  INV1S U26281 ( .I(gray_img[1975]), .O(n23150) );
  ND2S U26282 ( .I1(n20942), .I2(n23150), .O(n23159) );
  INV1S U26283 ( .I(n23159), .O(n20943) );
  NR2 U26284 ( .I1(gray_img[1983]), .I2(gray_img[1855]), .O(n23158) );
  AO12S U26285 ( .B1(n20943), .B2(n23158), .A1(n29680), .O(n20944) );
  ND2S U26286 ( .I1(n20945), .I2(n20944), .O(n13824) );
  AOI22S U26287 ( .A1(n25218), .A2(n25308), .B1(n25216), .B2(n25340), .O(
        n20946) );
  OA12S U26288 ( .B1(gray_img[647]), .B2(n29427), .A1(n29994), .O(n20947) );
  MOAI1S U26289 ( .A1(n29994), .A2(gray_img[647]), .B1(n25291), .B2(n20947), 
        .O(n20951) );
  INV1S U26290 ( .I(gray_img[1423]), .O(n20948) );
  INV1S U26291 ( .I(gray_img[1295]), .O(n29668) );
  ND2S U26292 ( .I1(n20948), .I2(n29668), .O(n29677) );
  INV1S U26293 ( .I(n29677), .O(n20949) );
  NR2 U26294 ( .I1(gray_img[1415]), .I2(gray_img[1287]), .O(n29676) );
  AO12S U26295 ( .B1(n20949), .B2(n29676), .A1(n29680), .O(n20950) );
  ND2S U26296 ( .I1(n20951), .I2(n20950), .O(n13978) );
  AOI22S U26297 ( .A1(n25086), .A2(n25162), .B1(n25085), .B2(n25361), .O(
        n20952) );
  OA12S U26298 ( .B1(gray_img[287]), .B2(n29427), .A1(n28248), .O(n20953) );
  MOAI1S U26299 ( .A1(n28248), .A2(gray_img[287]), .B1(n25291), .B2(n20953), 
        .O(n20957) );
  INV1S U26300 ( .I(gray_img[567]), .O(n20954) );
  INV1S U26301 ( .I(gray_img[695]), .O(n28169) );
  ND2S U26302 ( .I1(n20954), .I2(n28169), .O(n28178) );
  INV1S U26303 ( .I(n28178), .O(n20955) );
  NR2 U26304 ( .I1(gray_img[703]), .I2(gray_img[575]), .O(n28177) );
  AO12S U26305 ( .B1(n20955), .B2(n28177), .A1(n29680), .O(n20956) );
  ND2S U26306 ( .I1(n20957), .I2(n20956), .O(n13651) );
  AOI22S U26307 ( .A1(n25217), .A2(n25274), .B1(n25347), .B2(n25272), .O(
        n20958) );
  OA12S U26308 ( .B1(gray_img[919]), .B2(n29427), .A1(n30021), .O(n20959) );
  MOAI1S U26309 ( .A1(n30021), .A2(gray_img[919]), .B1(n25291), .B2(n20959), 
        .O(n20963) );
  INV1S U26310 ( .I(gray_img[1839]), .O(n20960) );
  ND2S U26311 ( .I1(n20960), .I2(n26681), .O(n26690) );
  INV1S U26312 ( .I(n26690), .O(n20961) );
  NR2 U26313 ( .I1(gray_img[1959]), .I2(gray_img[1831]), .O(n26689) );
  AO12S U26314 ( .B1(n20961), .B2(n26689), .A1(n29680), .O(n20962) );
  ND2S U26315 ( .I1(n20963), .I2(n20962), .O(n13828) );
  AOI22S U26316 ( .A1(n25326), .A2(n25273), .B1(n25325), .B2(n25271), .O(
        n20964) );
  OA12S U26317 ( .B1(gray_img[15]), .B2(n29427), .A1(n30081), .O(n20965) );
  MOAI1S U26318 ( .A1(n30081), .A2(gray_img[15]), .B1(n25291), .B2(n20965), 
        .O(n20969) );
  INV1S U26319 ( .I(gray_img[31]), .O(n20966) );
  INV1S U26320 ( .I(gray_img[159]), .O(n27876) );
  ND2S U26321 ( .I1(n20966), .I2(n27876), .O(n27885) );
  INV1S U26322 ( .I(n27885), .O(n20967) );
  NR2 U26323 ( .I1(gray_img[23]), .I2(gray_img[151]), .O(n27884) );
  AO12S U26324 ( .B1(n20967), .B2(n27884), .A1(n29680), .O(n20968) );
  ND2S U26325 ( .I1(n20969), .I2(n20968), .O(n13747) );
  AOI22S U26326 ( .A1(n25162), .A2(n25283), .B1(n25361), .B2(n25282), .O(
        n20970) );
  OA12S U26327 ( .B1(gray_img[319]), .B2(n29427), .A1(n26483), .O(n20971) );
  MOAI1S U26328 ( .A1(n26483), .A2(gray_img[319]), .B1(n25291), .B2(n20971), 
        .O(n20975) );
  INV1S U26329 ( .I(gray_img[631]), .O(n20972) );
  INV1S U26330 ( .I(gray_img[759]), .O(n26356) );
  ND2S U26331 ( .I1(n20972), .I2(n26356), .O(n26367) );
  INV1S U26332 ( .I(n26367), .O(n20973) );
  NR2 U26333 ( .I1(gray_img[767]), .I2(gray_img[639]), .O(n26366) );
  AO12S U26334 ( .B1(n20973), .B2(n26366), .A1(n29680), .O(n20974) );
  ND2S U26335 ( .I1(n20975), .I2(n20974), .O(n14135) );
  OA12S U26336 ( .B1(gray_img[47]), .B2(n29427), .A1(n26842), .O(n20976) );
  MOAI1S U26337 ( .A1(n26842), .A2(gray_img[47]), .B1(n25291), .B2(n20976), 
        .O(n20981) );
  INV1S U26338 ( .I(n20977), .O(n20979) );
  AO12S U26339 ( .B1(n20979), .B2(n20978), .A1(n29680), .O(n20980) );
  ND2S U26340 ( .I1(n20981), .I2(n20980), .O(n14241) );
  AOI22S U26341 ( .A1(n25308), .A2(n25245), .B1(n25340), .B2(n25244), .O(
        n20982) );
  OA12S U26342 ( .B1(gray_img[687]), .B2(n29427), .A1(n28601), .O(n20983) );
  MOAI1S U26343 ( .A1(n28601), .A2(gray_img[687]), .B1(n25291), .B2(n20983), 
        .O(n20987) );
  INV1S U26344 ( .I(gray_img[1503]), .O(n20984) );
  INV1S U26345 ( .I(gray_img[1375]), .O(n28372) );
  ND2S U26346 ( .I1(n20984), .I2(n28372), .O(n28393) );
  INV1S U26347 ( .I(n28393), .O(n20985) );
  NR2 U26348 ( .I1(gray_img[1367]), .I2(gray_img[1495]), .O(n28392) );
  AO12S U26349 ( .B1(n20985), .B2(n28392), .A1(n29680), .O(n20986) );
  ND2S U26350 ( .I1(n20987), .I2(n20986), .O(n13937) );
  AOI22S U26351 ( .A1(n25195), .A2(n25245), .B1(n25333), .B2(n25244), .O(
        n20988) );
  OA12S U26352 ( .B1(gray_img[559]), .B2(n29427), .A1(n28452), .O(n20989) );
  MOAI1S U26353 ( .A1(n28452), .A2(gray_img[559]), .B1(n25291), .B2(n20989), 
        .O(n20993) );
  INV1S U26354 ( .I(gray_img[1119]), .O(n20990) );
  INV1S U26355 ( .I(gray_img[1247]), .O(n28301) );
  ND2S U26356 ( .I1(n20990), .I2(n28301), .O(n28323) );
  INV1S U26357 ( .I(n28323), .O(n20991) );
  NR2 U26358 ( .I1(gray_img[1111]), .I2(gray_img[1239]), .O(n28322) );
  AO12S U26359 ( .B1(n20991), .B2(n28322), .A1(n29680), .O(n20992) );
  ND2S U26360 ( .I1(n20993), .I2(n20992), .O(n14021) );
  AOI22S U26361 ( .A1(n25086), .A2(n25195), .B1(n25085), .B2(n25333), .O(
        n20994) );
  OA12S U26362 ( .B1(gray_img[543]), .B2(n29427), .A1(n28943), .O(n20995) );
  MOAI1S U26363 ( .A1(n28943), .A2(gray_img[543]), .B1(n25291), .B2(n20995), 
        .O(n20999) );
  INV1S U26364 ( .I(gray_img[1087]), .O(n20996) );
  INV1S U26365 ( .I(gray_img[1215]), .O(n28865) );
  ND2S U26366 ( .I1(n20996), .I2(n28865), .O(n28887) );
  INV1S U26367 ( .I(n28887), .O(n20997) );
  NR2 U26368 ( .I1(gray_img[1207]), .I2(gray_img[1079]), .O(n28886) );
  AO12S U26369 ( .B1(n20997), .B2(n28886), .A1(n29680), .O(n20998) );
  ND2S U26370 ( .I1(n20999), .I2(n20998), .O(n14039) );
  AOI22S U26371 ( .A1(n25103), .A2(n25274), .B1(n25356), .B2(n25272), .O(
        n21000) );
  OA12S U26372 ( .B1(gray_img[791]), .B2(n29427), .A1(n29186), .O(n21001) );
  MOAI1S U26373 ( .A1(n29186), .A2(gray_img[791]), .B1(n25291), .B2(n21001), 
        .O(n21005) );
  INV1S U26374 ( .I(gray_img[1583]), .O(n21002) );
  INV1S U26375 ( .I(gray_img[1711]), .O(n29108) );
  ND2S U26376 ( .I1(n21002), .I2(n29108), .O(n29129) );
  INV1S U26377 ( .I(n29129), .O(n21003) );
  NR2 U26378 ( .I1(gray_img[1703]), .I2(gray_img[1575]), .O(n29128) );
  AO12S U26379 ( .B1(n21003), .B2(n29128), .A1(n29680), .O(n21004) );
  ND2S U26380 ( .I1(n21005), .I2(n21004), .O(n13890) );
  AOI22S U26381 ( .A1(n25162), .A2(n25326), .B1(n25361), .B2(n25325), .O(
        n21006) );
  OA12S U26382 ( .B1(gray_img[271]), .B2(n29427), .A1(n29374), .O(n21007) );
  MOAI1S U26383 ( .A1(n29374), .A2(gray_img[271]), .B1(n25291), .B2(n21007), 
        .O(n21011) );
  INV1S U26384 ( .I(gray_img[663]), .O(n21008) );
  ND2S U26385 ( .I1(n21008), .I2(n29062), .O(n29089) );
  INV1S U26386 ( .I(n29089), .O(n21009) );
  NR2 U26387 ( .I1(gray_img[671]), .I2(gray_img[543]), .O(n29088) );
  AO12S U26388 ( .B1(n21009), .B2(n29088), .A1(n29680), .O(n21010) );
  ND2S U26389 ( .I1(n21011), .I2(n21010), .O(n13700) );
  AOI22S U26390 ( .A1(n25372), .A2(n25283), .B1(n25370), .B2(n25282), .O(
        n21012) );
  OA12S U26391 ( .B1(gray_img[447]), .B2(n29427), .A1(n26466), .O(n21013) );
  MOAI1S U26392 ( .A1(n26466), .A2(gray_img[447]), .B1(n25291), .B2(n21013), 
        .O(n21017) );
  INV1S U26393 ( .I(gray_img[1015]), .O(n21014) );
  ND2S U26394 ( .I1(n21014), .I2(n26387), .O(n26409) );
  INV1S U26395 ( .I(n26409), .O(n21015) );
  NR2 U26396 ( .I1(gray_img[895]), .I2(gray_img[1023]), .O(n26408) );
  AO12S U26397 ( .B1(n21015), .B2(n26408), .A1(n29680), .O(n21016) );
  ND2S U26398 ( .I1(n21017), .I2(n21016), .O(n14091) );
  AOI22S U26399 ( .A1(n25218), .A2(n25162), .B1(n25216), .B2(n25361), .O(
        n21018) );
  OA12S U26400 ( .B1(gray_img[263]), .B2(n29427), .A1(n30006), .O(n21019) );
  MOAI1S U26401 ( .A1(n30006), .A2(gray_img[263]), .B1(n25291), .B2(n21019), 
        .O(n21022) );
  INV1S U26402 ( .I(gray_img[527]), .O(n25136) );
  INV1S U26403 ( .I(gray_img[655]), .O(n29917) );
  ND2S U26404 ( .I1(n25136), .I2(n29917), .O(n29938) );
  INV1S U26405 ( .I(n29938), .O(n21020) );
  NR2 U26406 ( .I1(gray_img[519]), .I2(gray_img[647]), .O(n29937) );
  AO12S U26407 ( .B1(n21020), .B2(n29937), .A1(n29680), .O(n21021) );
  ND2S U26408 ( .I1(n21022), .I2(n21021), .O(n13729) );
  AOI22S U26409 ( .A1(n25246), .A2(n25283), .B1(n25257), .B2(n25282), .O(
        n21023) );
  OA12S U26410 ( .B1(gray_img[191]), .B2(n29427), .A1(n27685), .O(n21024) );
  MOAI1S U26411 ( .A1(n27685), .A2(gray_img[191]), .B1(n25291), .B2(n21024), 
        .O(n21028) );
  INV1S U26412 ( .I(gray_img[383]), .O(n21025) );
  INV1S U26413 ( .I(gray_img[511]), .O(n27622) );
  ND2S U26414 ( .I1(n21025), .I2(n27622), .O(n27629) );
  INV1S U26415 ( .I(n27629), .O(n21026) );
  NR2 U26416 ( .I1(gray_img[503]), .I2(gray_img[375]), .O(n27628) );
  AO12S U26417 ( .B1(n21026), .B2(n27628), .A1(n29680), .O(n21027) );
  ND2S U26418 ( .I1(n21028), .I2(n21027), .O(n14179) );
  AOI22S U26419 ( .A1(n25373), .A2(n25246), .B1(n25371), .B2(n25257), .O(
        n21029) );
  OA12S U26420 ( .B1(gray_img[183]), .B2(n29427), .A1(n27779), .O(n21030) );
  MOAI1S U26421 ( .A1(n27779), .A2(gray_img[183]), .B1(n25291), .B2(n21030), 
        .O(n21034) );
  INV1S U26422 ( .I(gray_img[495]), .O(n21031) );
  INV1S U26423 ( .I(gray_img[367]), .O(n27463) );
  ND2S U26424 ( .I1(n21031), .I2(n27463), .O(n27484) );
  INV1S U26425 ( .I(n27484), .O(n21032) );
  NR2 U26426 ( .I1(gray_img[487]), .I2(gray_img[359]), .O(n27483) );
  AO12S U26427 ( .B1(n21032), .B2(n27483), .A1(n29680), .O(n21033) );
  ND2S U26428 ( .I1(n21034), .I2(n21033), .O(n14188) );
  AOI22S U26429 ( .A1(n25373), .A2(n25195), .B1(n25371), .B2(n25333), .O(
        n21035) );
  OA12S U26430 ( .B1(gray_img[567]), .B2(n29427), .A1(n28121), .O(n21036) );
  MOAI1S U26431 ( .A1(n28121), .A2(gray_img[567]), .B1(n25291), .B2(n21036), 
        .O(n21040) );
  INV1S U26432 ( .I(gray_img[1263]), .O(n21037) );
  INV1S U26433 ( .I(gray_img[1135]), .O(n28055) );
  ND2S U26434 ( .I1(n21037), .I2(n28055), .O(n28062) );
  INV1S U26435 ( .I(n28062), .O(n21038) );
  NR2 U26436 ( .I1(gray_img[1255]), .I2(gray_img[1127]), .O(n28061) );
  AO12S U26437 ( .B1(n21038), .B2(n28061), .A1(n29680), .O(n21039) );
  ND2S U26438 ( .I1(n21040), .I2(n21039), .O(n14012) );
  AOI22S U26439 ( .A1(n25273), .A2(n25283), .B1(n25271), .B2(n25282), .O(
        n21041) );
  OA12S U26440 ( .B1(gray_img[63]), .B2(n29427), .A1(n27702), .O(n21042) );
  MOAI1S U26441 ( .A1(n27702), .A2(gray_img[63]), .B1(n25291), .B2(n21042), 
        .O(n21046) );
  INV1S U26442 ( .I(gray_img[119]), .O(n21043) );
  INV1S U26443 ( .I(gray_img[247]), .O(n27580) );
  ND2S U26444 ( .I1(n21043), .I2(n27580), .O(n27591) );
  INV1S U26445 ( .I(n27591), .O(n21044) );
  NR2 U26446 ( .I1(gray_img[255]), .I2(gray_img[127]), .O(n27590) );
  AO12S U26447 ( .B1(n21044), .B2(n27590), .A1(n29680), .O(n21045) );
  ND2S U26448 ( .I1(n21046), .I2(n21045), .O(n14223) );
  AOI22S U26449 ( .A1(n25373), .A2(n25308), .B1(n25371), .B2(n25340), .O(
        n21047) );
  OA12S U26450 ( .B1(gray_img[695]), .B2(n29427), .A1(n28208), .O(n21048) );
  MOAI1S U26451 ( .A1(n28208), .A2(gray_img[695]), .B1(n25291), .B2(n21048), 
        .O(n21052) );
  INV1S U26452 ( .I(gray_img[1391]), .O(n21049) );
  INV1S U26453 ( .I(gray_img[1519]), .O(n27984) );
  ND2S U26454 ( .I1(n21049), .I2(n27984), .O(n28011) );
  INV1S U26455 ( .I(n28011), .O(n21050) );
  NR2 U26456 ( .I1(gray_img[1383]), .I2(gray_img[1511]), .O(n28010) );
  AO12S U26457 ( .B1(n21050), .B2(n28010), .A1(n29680), .O(n21051) );
  ND2S U26458 ( .I1(n21052), .I2(n21051), .O(n13930) );
  AOI22S U26459 ( .A1(n25086), .A2(n25273), .B1(n25085), .B2(n25271), .O(
        n21053) );
  OA12S U26460 ( .B1(gray_img[31]), .B2(n29427), .A1(n27814), .O(n21054) );
  MOAI1S U26461 ( .A1(n27814), .A2(gray_img[31]), .B1(n25291), .B2(n21054), 
        .O(n21058) );
  INV1S U26462 ( .I(gray_img[191]), .O(n21055) );
  INV1S U26463 ( .I(gray_img[63]), .O(n27721) );
  ND2S U26464 ( .I1(n21055), .I2(n27721), .O(n27743) );
  INV1S U26465 ( .I(n27743), .O(n21056) );
  NR2 U26466 ( .I1(gray_img[55]), .I2(gray_img[183]), .O(n27742) );
  AO12S U26467 ( .B1(n21056), .B2(n27742), .A1(n29680), .O(n21057) );
  ND2S U26468 ( .I1(n21058), .I2(n21057), .O(n13785) );
  AOI22S U26469 ( .A1(n25308), .A2(n25274), .B1(n25340), .B2(n25272), .O(
        n21059) );
  OA12S U26470 ( .B1(gray_img[663]), .B2(n29427), .A1(n29033), .O(n21060) );
  MOAI1S U26471 ( .A1(n29033), .A2(gray_img[663]), .B1(n25291), .B2(n21060), 
        .O(n21064) );
  INV1S U26472 ( .I(gray_img[1327]), .O(n21061) );
  INV1S U26473 ( .I(gray_img[1455]), .O(n28974) );
  ND2S U26474 ( .I1(n21061), .I2(n28974), .O(n28981) );
  INV1S U26475 ( .I(n28981), .O(n21062) );
  NR2 U26476 ( .I1(gray_img[1447]), .I2(gray_img[1319]), .O(n28980) );
  AO12S U26477 ( .B1(n21062), .B2(n28980), .A1(n29680), .O(n21063) );
  ND2S U26478 ( .I1(n21064), .I2(n21063), .O(n13960) );
  AOI22S U26479 ( .A1(n25217), .A2(n25283), .B1(n25347), .B2(n25282), .O(
        n21065) );
  OA12S U26480 ( .B1(gray_img[959]), .B2(n29427), .A1(n28718), .O(n21066) );
  MOAI1S U26481 ( .A1(n28718), .A2(gray_img[959]), .B1(n25291), .B2(n21066), 
        .O(n21070) );
  INV1S U26482 ( .I(gray_img[1911]), .O(n21067) );
  INV1S U26483 ( .I(gray_img[2039]), .O(n25969) );
  ND2S U26484 ( .I1(n21067), .I2(n25969), .O(n25976) );
  INV1S U26485 ( .I(n25976), .O(n21068) );
  NR2 U26486 ( .I1(gray_img[2047]), .I2(gray_img[1919]), .O(n25975) );
  AO12S U26487 ( .B1(n21068), .B2(n25975), .A1(n29680), .O(n21069) );
  ND2S U26488 ( .I1(n21070), .I2(n21069), .O(n15468) );
  AOI22S U26489 ( .A1(n25246), .A2(n25274), .B1(n25257), .B2(n25272), .O(
        n21071) );
  OA12S U26490 ( .B1(gray_img[151]), .B2(n29427), .A1(n30070), .O(n21072) );
  MOAI1S U26491 ( .A1(n30070), .A2(gray_img[151]), .B1(n25291), .B2(n21072), 
        .O(n21076) );
  INV1S U26492 ( .I(gray_img[423]), .O(n21073) );
  INV1S U26493 ( .I(gray_img[295]), .O(n27275) );
  ND2S U26494 ( .I1(n21073), .I2(n27275), .O(n27296) );
  INV1S U26495 ( .I(n27296), .O(n21074) );
  NR2 U26496 ( .I1(gray_img[303]), .I2(gray_img[431]), .O(n27295) );
  AO12S U26497 ( .B1(n21074), .B2(n27295), .A1(n29680), .O(n21075) );
  ND2S U26498 ( .I1(n21076), .I2(n21075), .O(n13765) );
  AOI22S U26499 ( .A1(n25373), .A2(n25103), .B1(n25371), .B2(n25356), .O(
        n21077) );
  OA12S U26500 ( .B1(gray_img[823]), .B2(n29427), .A1(n25929), .O(n21078) );
  MOAI1S U26501 ( .A1(n25929), .A2(gray_img[823]), .B1(n25291), .B2(n21078), 
        .O(n21082) );
  INV1S U26502 ( .I(gray_img[1775]), .O(n21079) );
  ND2S U26503 ( .I1(n21079), .I2(n25792), .O(n25813) );
  INV1S U26504 ( .I(n25813), .O(n21080) );
  NR2 U26505 ( .I1(gray_img[1639]), .I2(gray_img[1767]), .O(n25812) );
  AO12S U26506 ( .B1(n21080), .B2(n25812), .A1(n29680), .O(n21081) );
  ND2S U26507 ( .I1(n21082), .I2(n21081), .O(n13866) );
  AOI22S U26508 ( .A1(n25103), .A2(n25086), .B1(n25356), .B2(n25085), .O(
        n21083) );
  OA12S U26509 ( .B1(gray_img[799]), .B2(n29427), .A1(n29266), .O(n21084) );
  MOAI1S U26510 ( .A1(n29266), .A2(gray_img[799]), .B1(n25291), .B2(n21084), 
        .O(n21088) );
  INV1S U26511 ( .I(gray_img[1591]), .O(n21085) );
  INV1S U26512 ( .I(gray_img[1719]), .O(n29221) );
  ND2S U26513 ( .I1(n21085), .I2(n29221), .O(n29230) );
  INV1S U26514 ( .I(n29230), .O(n21086) );
  NR2 U26515 ( .I1(gray_img[1727]), .I2(gray_img[1599]), .O(n29229) );
  AO12S U26516 ( .B1(n21086), .B2(n29229), .A1(n29680), .O(n21087) );
  ND2S U26517 ( .I1(n21088), .I2(n21087), .O(n13884) );
  NR2 U26518 ( .I1(cnt_dyn[2]), .I2(n30307), .O(n22782) );
  INV1S U26519 ( .I(n30251), .O(n30424) );
  AOI22S U26520 ( .A1(n21089), .A2(gray_img[222]), .B1(gray_img[1246]), .B2(
        n21090), .O(n21095) );
  NR2 U26521 ( .I1(cnt_bdyn[0]), .I2(n30369), .O(n30135) );
  NR2 U26522 ( .I1(n21151), .I2(n21146), .O(n22735) );
  INV1S U26523 ( .I(n22735), .O(n22884) );
  INV1S U26524 ( .I(n22884), .O(n22785) );
  AOI22S U26525 ( .A1(n22785), .A2(gray_img[350]), .B1(gray_img[838]), .B2(
        n22513), .O(n21094) );
  NR2 U26526 ( .I1(n21158), .I2(n21144), .O(n22896) );
  INV1S U26527 ( .I(n22540), .O(n22796) );
  ND2S U26528 ( .I1(n22796), .I2(gray_img[1750]), .O(n21093) );
  NR2 U26529 ( .I1(n21151), .I2(n21147), .O(n22867) );
  INV1S U26530 ( .I(n22867), .O(n22725) );
  INV1S U26531 ( .I(gray_img[862]), .O(n23076) );
  NR2 U26532 ( .I1(cnt_dyn[1]), .I2(n30333), .O(n30298) );
  INV1S U26533 ( .I(n22865), .O(n22837) );
  AOI22S U26534 ( .A1(n22837), .A2(gray_img[334]), .B1(gray_img[1118]), .B2(
        n22935), .O(n21091) );
  OAI12HS U26535 ( .B1(n22725), .B2(n23076), .A1(n21091), .O(n21092) );
  AN4B1S U26536 ( .I1(n21095), .I2(n21094), .I3(n21093), .B1(n21092), .O(
        n21171) );
  NR2 U26537 ( .I1(n30364), .I2(n21138), .O(n22828) );
  NR2 U26538 ( .I1(n21153), .I2(n21144), .O(n22827) );
  AOI22S U26539 ( .A1(n22828), .A2(gray_img[982]), .B1(gray_img[1622]), .B2(
        n15919), .O(n21102) );
  NR2 U26540 ( .I1(n21154), .I2(n21147), .O(n22787) );
  INV1S U26541 ( .I(n22787), .O(n21504) );
  INV1S U26542 ( .I(n21504), .O(n22864) );
  NR2 U26543 ( .I1(n21145), .I2(n21147), .O(n22794) );
  AOI22S U26544 ( .A1(n22864), .A2(gray_img[1886]), .B1(gray_img[1862]), .B2(
        n22794), .O(n21101) );
  ND2S U26545 ( .I1(n21096), .I2(gray_img[1502]), .O(n21100) );
  NR2 U26546 ( .I1(n21156), .I2(n21144), .O(n22809) );
  INV1S U26547 ( .I(n15921), .O(n22058) );
  INV1S U26548 ( .I(n21097), .O(n22670) );
  INV1S U26549 ( .I(gray_img[1606]), .O(n25676) );
  MOAI1S U26550 ( .A1(n22670), .A2(n25676), .B1(gray_img[214]), .B2(n15918), 
        .O(n21098) );
  AO12S U26551 ( .B1(gray_img[1238]), .B2(n15921), .A1(n21098), .O(n21099) );
  AN4B1S U26552 ( .I1(n21102), .I2(n21101), .I3(n21100), .B1(n21099), .O(
        n21170) );
  NR2 U26553 ( .I1(n21144), .I2(n21146), .O(n22889) );
  AOI22S U26554 ( .A1(n22863), .A2(gray_img[1878]), .B1(gray_img[1366]), .B2(
        n22889), .O(n21105) );
  NR2 U26555 ( .I1(n30364), .I2(n21131), .O(n22911) );
  AOI22S U26556 ( .A1(n22911), .A2(gray_img[966]), .B1(gray_img[454]), .B2(
        n22686), .O(n21104) );
  NR2 U26557 ( .I1(n30364), .I2(n21114), .O(n22910) );
  NR2 U26558 ( .I1(n21158), .I2(n21114), .O(n22888) );
  AOI22S U26559 ( .A1(n22910), .A2(gray_img[974]), .B1(gray_img[718]), .B2(
        n22888), .O(n21103) );
  ND3S U26560 ( .I1(n21105), .I2(n21104), .I3(n21103), .O(n21113) );
  NR2 U26561 ( .I1(n21156), .I2(n21145), .O(n22838) );
  INV1S U26562 ( .I(n22838), .O(n22392) );
  INV1S U26563 ( .I(gray_img[1222]), .O(n28504) );
  MOAI1S U26564 ( .A1(n22392), .A2(n28504), .B1(n22770), .B2(gray_img[1734]), 
        .O(n21108) );
  INV1S U26565 ( .I(n21106), .O(n22718) );
  INV1S U26566 ( .I(gray_img[1478]), .O(n23510) );
  MOAI1S U26567 ( .A1(n22718), .A2(n23510), .B1(n22625), .B2(gray_img[326]), 
        .O(n21107) );
  NR2 U26568 ( .I1(n21108), .I2(n21107), .O(n21111) );
  NR2 U26569 ( .I1(n21153), .I2(n21114), .O(n22887) );
  NR2 U26570 ( .I1(n21158), .I2(n21154), .O(n22505) );
  AOI22S U26571 ( .A1(n22887), .A2(gray_img[590]), .B1(gray_img[1758]), .B2(
        n22505), .O(n21110) );
  INV1S U26572 ( .I(n22803), .O(n22883) );
  NR2 U26573 ( .I1(n21151), .I2(n21157), .O(n22736) );
  AOI22S U26574 ( .A1(n22883), .A2(gray_img[734]), .B1(gray_img[478]), .B2(
        n22736), .O(n21109) );
  ND3S U26575 ( .I1(n21111), .I2(n21110), .I3(n21109), .O(n21112) );
  NR2 U26576 ( .I1(n21113), .I2(n21112), .O(n21168) );
  NR2 U26577 ( .I1(n23571), .I2(n22853), .O(n21119) );
  NR2 U26578 ( .I1(n21153), .I2(n21138), .O(n22945) );
  ND2S U26579 ( .I1(n15915), .I2(gray_img[598]), .O(n21117) );
  NR2 U26580 ( .I1(n21114), .I2(n21147), .O(n22724) );
  BUF1 U26581 ( .I(n22724), .O(n22932) );
  AOI22S U26582 ( .A1(n22610), .A2(gray_img[198]), .B1(gray_img[846]), .B2(
        n22932), .O(n21116) );
  NR2 U26583 ( .I1(n21114), .I2(n21156), .O(n22836) );
  NR2 U26584 ( .I1(n21114), .I2(n21157), .O(n22862) );
  AOI22S U26585 ( .A1(n22836), .A2(gray_img[206]), .B1(gray_img[462]), .B2(
        n22862), .O(n21115) );
  ND3S U26586 ( .I1(n21117), .I2(n21116), .I3(n21115), .O(n21118) );
  NR2 U26587 ( .I1(n21119), .I2(n21118), .O(n21167) );
  ND2S U26588 ( .I1(n22893), .I2(gray_img[70]), .O(n21136) );
  NR2 U26589 ( .I1(n21158), .I2(n21138), .O(n22920) );
  INV1S U26590 ( .I(n22920), .O(n21933) );
  AOI22S U26591 ( .A1(n22695), .A2(gray_img[726]), .B1(gray_img[1494]), .B2(
        n22664), .O(n21135) );
  NR2 U26592 ( .I1(n30364), .I2(n21151), .O(n22873) );
  INV1S U26593 ( .I(n22873), .O(n22682) );
  INV1S U26594 ( .I(n22682), .O(n22819) );
  ND2S U26595 ( .I1(n22819), .I2(gray_img[990]), .O(n21130) );
  NR2 U26596 ( .I1(n21147), .I2(n21138), .O(n21121) );
  BUF1 U26597 ( .I(n21121), .O(n22930) );
  AOI22S U26598 ( .A1(gray_img[1374]), .A2(n21120), .B1(gray_img[854]), .B2(
        n22930), .O(n21124) );
  AOI22S U26599 ( .A1(gray_img[2006]), .A2(n22679), .B1(gray_img[342]), .B2(
        n15905), .O(n21123) );
  AN2 U26600 ( .I1(n30451), .I2(n30322), .O(n22901) );
  ND2S U26601 ( .I1(gray_img[86]), .I2(n22901), .O(n21122) );
  ND3S U26602 ( .I1(n21124), .I2(n21123), .I3(n21122), .O(n21128) );
  NR2 U26603 ( .I1(n23599), .I2(n22811), .O(n21127) );
  AN2 U26604 ( .I1(n30299), .I2(n21125), .O(n22812) );
  INV1S U26605 ( .I(n22812), .O(n22904) );
  NR2 U26606 ( .I1(n23558), .I2(n22904), .O(n21126) );
  NR3 U26607 ( .I1(n21128), .I2(n21127), .I3(n21126), .O(n21129) );
  ND2S U26608 ( .I1(n21130), .I2(n21129), .O(n21133) );
  NR2 U26609 ( .I1(n21158), .I2(n21131), .O(n22909) );
  INV1S U26610 ( .I(n22909), .O(n22156) );
  MOAI1S U26611 ( .A1(n22156), .A2(n27144), .B1(n22630), .B2(gray_img[582]), 
        .O(n21132) );
  NR2 U26612 ( .I1(n21133), .I2(n21132), .O(n21134) );
  ND3S U26613 ( .I1(n21136), .I2(n21135), .I3(n21134), .O(n21143) );
  INV1S U26614 ( .I(n30322), .O(n30308) );
  INV1S U26615 ( .I(n21137), .O(n22924) );
  NR2 U26616 ( .I1(n30251), .I2(n30361), .O(n22755) );
  INV1S U26617 ( .I(n22755), .O(n22251) );
  INV1S U26618 ( .I(n22251), .O(n22919) );
  ND2S U26619 ( .I1(n22919), .I2(gray_img[2014]), .O(n21140) );
  NR2 U26620 ( .I1(n21159), .I2(n21153), .O(n22656) );
  NR2 U26621 ( .I1(n21157), .I2(n21138), .O(n22895) );
  AOI22S U26622 ( .A1(n22656), .A2(gray_img[1614]), .B1(n22895), .B2(
        gray_img[470]), .O(n21139) );
  OAI112HS U26623 ( .C1(n22924), .C2(n21141), .A1(n21140), .B1(n21139), .O(
        n21142) );
  NR2 U26624 ( .I1(n21143), .I2(n21142), .O(n21166) );
  NR2 U26625 ( .I1(n30306), .I2(n21144), .O(n22663) );
  INV1S U26626 ( .I(n22663), .O(n21842) );
  INV1S U26627 ( .I(n21842), .O(n22929) );
  ND2S U26628 ( .I1(n22929), .I2(gray_img[1110]), .O(n21150) );
  AOI22S U26629 ( .A1(n22934), .A2(gray_img[1350]), .B1(gray_img[1094]), .B2(
        n22703), .O(n21149) );
  NR2 U26630 ( .I1(n21159), .I2(n21146), .O(n22846) );
  NR2 U26631 ( .I1(n21159), .I2(n21147), .O(n22937) );
  AOI22S U26632 ( .A1(n22846), .A2(gray_img[1358]), .B1(gray_img[1870]), .B2(
        n22937), .O(n21148) );
  ND3S U26633 ( .I1(n21150), .I2(n21149), .I3(n21148), .O(n21164) );
  NR2 U26634 ( .I1(n21154), .I2(n21153), .O(n22694) );
  AOI22S U26635 ( .A1(n21152), .A2(gray_img[606]), .B1(gray_img[1630]), .B2(
        n22694), .O(n21162) );
  AOI22S U26636 ( .A1(n21155), .A2(gray_img[1102]), .B1(gray_img[1230]), .B2(
        n22936), .O(n21161) );
  NR2 U26637 ( .I1(n21159), .I2(n21157), .O(n22369) );
  INV1S U26638 ( .I(n22487), .O(n22921) );
  AOI22S U26639 ( .A1(n22369), .A2(gray_img[1486]), .B1(gray_img[1742]), .B2(
        n22921), .O(n21160) );
  ND3S U26640 ( .I1(n21162), .I2(n21161), .I3(n21160), .O(n21163) );
  NR2 U26641 ( .I1(n21164), .I2(n21163), .O(n21165) );
  AN4S U26642 ( .I1(n21168), .I2(n21167), .I3(n21166), .I4(n21165), .O(n21169)
         );
  ND3S U26643 ( .I1(n21171), .I2(n21170), .I3(n21169), .O(n21224) );
  NR2 U26644 ( .I1(cnt_dyn[3]), .I2(n30305), .O(n22957) );
  INV1S U26645 ( .I(n15919), .O(n22601) );
  AOI22S U26646 ( .A1(n21155), .A2(gray_img[1070]), .B1(n22827), .B2(
        gray_img[1590]), .O(n21175) );
  AOI22S U26647 ( .A1(n22810), .A2(gray_img[678]), .B1(gray_img[558]), .B2(
        n22887), .O(n21174) );
  BUF1 U26648 ( .I(n22862), .O(n22762) );
  AOI22S U26649 ( .A1(n22625), .A2(gray_img[294]), .B1(gray_img[430]), .B2(
        n22762), .O(n21173) );
  INV1S U26650 ( .I(gray_img[1446]), .O(n28960) );
  MOAI1S U26651 ( .A1(n22718), .A2(n28960), .B1(n22838), .B2(gray_img[1190]), 
        .O(n21172) );
  AN4B1S U26652 ( .I1(n21175), .I2(n21174), .I3(n21173), .B1(n21172), .O(
        n21222) );
  AOI22S U26653 ( .A1(n22828), .A2(gray_img[950]), .B1(gray_img[1462]), .B2(
        n22664), .O(n21181) );
  AOI22S U26654 ( .A1(n22864), .A2(gray_img[1854]), .B1(gray_img[1198]), .B2(
        n22936), .O(n21180) );
  ND2S U26655 ( .I1(n22863), .I2(gray_img[1846]), .O(n21179) );
  ND2S U26656 ( .I1(n22889), .I2(gray_img[1334]), .O(n21177) );
  AOI22S U26657 ( .A1(gray_img[1342]), .A2(n21120), .B1(n22630), .B2(
        gray_img[550]), .O(n21176) );
  ND2S U26658 ( .I1(n21177), .I2(n21176), .O(n21178) );
  AN4B1S U26659 ( .I1(n21181), .I2(n21180), .I3(n21179), .B1(n21178), .O(
        n21221) );
  NR2 U26660 ( .I1(n26679), .I2(n22853), .O(n21194) );
  ND2S U26661 ( .I1(n22929), .I2(gray_img[1078]), .O(n21184) );
  AOI22S U26662 ( .A1(n22837), .A2(gray_img[302]), .B1(gray_img[1086]), .B2(
        n22935), .O(n21183) );
  INV1S U26663 ( .I(n22794), .O(n22364) );
  INV1S U26664 ( .I(n22364), .O(n22938) );
  AOI22S U26665 ( .A1(n22938), .A2(gray_img[1830]), .B1(gray_img[1062]), .B2(
        n22703), .O(n21182) );
  ND3S U26666 ( .I1(n21184), .I2(n21183), .I3(n21182), .O(n21193) );
  ND2S U26667 ( .I1(n21152), .I2(gray_img[574]), .O(n21188) );
  INV1S U26668 ( .I(n22846), .O(n22031) );
  INV1S U26669 ( .I(n22031), .O(n22861) );
  AOI22S U26670 ( .A1(n22861), .A2(gray_img[1326]), .B1(gray_img[1838]), .B2(
        n22937), .O(n21187) );
  INV1S U26671 ( .I(n22369), .O(n22875) );
  INV1S U26672 ( .I(n22875), .O(n22847) );
  AOI22S U26673 ( .A1(n22934), .A2(gray_img[1318]), .B1(gray_img[1454]), .B2(
        n22847), .O(n21186) );
  INV1S U26674 ( .I(gray_img[1710]), .O(n29106) );
  MOAI1S U26675 ( .A1(n22487), .A2(n29106), .B1(n22656), .B2(gray_img[1582]), 
        .O(n21185) );
  AN4B1S U26676 ( .I1(n21188), .I2(n21187), .I3(n21186), .B1(n21185), .O(
        n21191) );
  AOI22S U26677 ( .A1(n22867), .A2(gray_img[830]), .B1(gray_img[190]), .B2(
        n21089), .O(n21190) );
  AOI22S U26678 ( .A1(n21096), .A2(gray_img[1470]), .B1(gray_img[1598]), .B2(
        n22694), .O(n21189) );
  NR3 U26679 ( .I1(n21194), .I2(n21193), .I3(n21192), .O(n21219) );
  ND2S U26680 ( .I1(n15918), .I2(gray_img[182]), .O(n21206) );
  AOI22S U26681 ( .A1(n22883), .A2(gray_img[702]), .B1(gray_img[318]), .B2(
        n22735), .O(n21205) );
  AOI22S U26682 ( .A1(n22770), .A2(gray_img[1702]), .B1(gray_img[1574]), .B2(
        n21097), .O(n21204) );
  INV1S U26683 ( .I(gray_img[46]), .O(n26966) );
  AOI22S U26684 ( .A1(gray_img[54]), .A2(n22901), .B1(gray_img[1974]), .B2(
        n22679), .O(n21196) );
  ND2S U26685 ( .I1(n22812), .I2(gray_img[1958]), .O(n21195) );
  OAI112HS U26686 ( .C1(n22811), .C2(n26966), .A1(n21196), .B1(n21195), .O(
        n21199) );
  INV1S U26687 ( .I(gray_img[958]), .O(n26121) );
  NR2 U26688 ( .I1(n26121), .I2(n22682), .O(n21198) );
  INV1S U26689 ( .I(n22911), .O(n21841) );
  INV1S U26690 ( .I(gray_img[934]), .O(n23230) );
  MOAI1S U26691 ( .A1(n21841), .A2(n23230), .B1(n22686), .B2(gray_img[422]), 
        .O(n21197) );
  NR3 U26692 ( .I1(n21199), .I2(n21198), .I3(n21197), .O(n21202) );
  INV1S U26693 ( .I(n22910), .O(n22346) );
  AOI22S U26694 ( .A1(n22802), .A2(gray_img[942]), .B1(gray_img[686]), .B2(
        n22888), .O(n21201) );
  INV1S U26695 ( .I(n22505), .O(n22882) );
  INV1S U26696 ( .I(n22882), .O(n22786) );
  AOI22S U26697 ( .A1(n22786), .A2(gray_img[1726]), .B1(gray_img[446]), .B2(
        n22736), .O(n21200) );
  ND3S U26698 ( .I1(n21202), .I2(n21201), .I3(n21200), .O(n21203) );
  AN4B1S U26699 ( .I1(n21206), .I2(n21205), .I3(n21204), .B1(n21203), .O(
        n21218) );
  AOI22S U26700 ( .A1(n22513), .A2(gray_img[806]), .B1(gray_img[166]), .B2(
        n22610), .O(n21210) );
  AOI22S U26701 ( .A1(n22836), .A2(gray_img[174]), .B1(gray_img[814]), .B2(
        n22932), .O(n21209) );
  ND2S U26702 ( .I1(n15905), .I2(gray_img[310]), .O(n21208) );
  INV1S U26703 ( .I(n22930), .O(n22841) );
  INV1S U26704 ( .I(gray_img[822]), .O(n26108) );
  MOAI1S U26705 ( .A1(n22841), .A2(n26108), .B1(n15915), .B2(gray_img[566]), 
        .O(n21207) );
  AN4B1S U26706 ( .I1(n21210), .I2(n21209), .I3(n21208), .B1(n21207), .O(
        n21217) );
  ND2S U26707 ( .I1(n22893), .I2(gray_img[38]), .O(n21213) );
  AOI22S U26708 ( .A1(n22895), .A2(gray_img[438]), .B1(gray_img[694]), .B2(
        n22920), .O(n21212) );
  AOI22S U26709 ( .A1(n22896), .A2(gray_img[1718]), .B1(gray_img[1206]), .B2(
        n15921), .O(n21211) );
  ND3S U26710 ( .I1(n21213), .I2(n21212), .I3(n21211), .O(n21215) );
  MOAI1S U26711 ( .A1(n22924), .A2(n27719), .B1(gray_img[1214]), .B2(n21090), 
        .O(n21214) );
  AO112S U26712 ( .C1(gray_img[1982]), .C2(n22919), .A1(n21215), .B1(n21214), 
        .O(n21216) );
  AN4B1S U26713 ( .I1(n21219), .I2(n21218), .I3(n21217), .B1(n21216), .O(
        n21220) );
  ND3S U26714 ( .I1(n21222), .I2(n21221), .I3(n21220), .O(n21223) );
  AOI22S U26715 ( .A1(n22782), .A2(n21224), .B1(n22957), .B2(n21223), .O(
        n21336) );
  INV1S U26716 ( .I(n30281), .O(n22784) );
  MOAI1S U26717 ( .A1(n22392), .A2(n26637), .B1(n22610), .B2(gray_img[134]), 
        .O(n21230) );
  MOAI1S U26718 ( .A1(n22865), .A2(n21225), .B1(n22836), .B2(gray_img[142]), 
        .O(n21229) );
  INV1S U26719 ( .I(n21152), .O(n22750) );
  AOI22S U26720 ( .A1(n22630), .A2(gray_img[518]), .B1(gray_img[902]), .B2(
        n22566), .O(n21227) );
  ND2S U26721 ( .I1(n22695), .I2(gray_img[662]), .O(n21226) );
  OAI112HS U26722 ( .C1(n22750), .C2(n29076), .A1(n21227), .B1(n21226), .O(
        n21228) );
  NR3 U26723 ( .I1(n21230), .I2(n21229), .I3(n21228), .O(n21276) );
  INV1S U26724 ( .I(gray_img[1414]), .O(n29654) );
  MOAI1S U26725 ( .A1(n22718), .A2(n29654), .B1(n22883), .B2(gray_img[670]), 
        .O(n21235) );
  INV1S U26726 ( .I(n22895), .O(n22658) );
  INV1S U26727 ( .I(gray_img[406]), .O(n28744) );
  MOAI1S U26728 ( .A1(n22658), .A2(n28744), .B1(gray_img[1030]), .B2(n22703), 
        .O(n21234) );
  INV1S U26729 ( .I(gray_img[1686]), .O(n26556) );
  ND2S U26730 ( .I1(n15915), .I2(gray_img[534]), .O(n21232) );
  INV1S U26731 ( .I(n22736), .O(n21288) );
  INV1S U26732 ( .I(n21288), .O(n22881) );
  AOI22S U26733 ( .A1(gray_img[158]), .A2(n21089), .B1(n22881), .B2(
        gray_img[414]), .O(n21231) );
  OAI112HS U26734 ( .C1(n22540), .C2(n26556), .A1(n21232), .B1(n21231), .O(
        n21233) );
  NR3 U26735 ( .I1(n21235), .I2(n21234), .I3(n21233), .O(n21275) );
  INV1S U26736 ( .I(gray_img[1950]), .O(n29514) );
  AOI22S U26737 ( .A1(n22369), .A2(gray_img[1422]), .B1(gray_img[1678]), .B2(
        n22921), .O(n21239) );
  INV1S U26738 ( .I(n22725), .O(n22813) );
  ND2S U26739 ( .I1(n22813), .I2(gray_img[798]), .O(n21238) );
  AOI22S U26740 ( .A1(n22656), .A2(gray_img[1550]), .B1(gray_img[1294]), .B2(
        n22846), .O(n21237) );
  INV1S U26741 ( .I(n21155), .O(n22848) );
  INV1S U26742 ( .I(gray_img[1038]), .O(n26625) );
  MOAI1S U26743 ( .A1(n22848), .A2(n26625), .B1(n22936), .B2(gray_img[1166]), 
        .O(n21236) );
  AN4B1S U26744 ( .I1(n21239), .I2(n21238), .I3(n21237), .B1(n21236), .O(
        n21241) );
  AOI22S U26745 ( .A1(n21096), .A2(gray_img[1438]), .B1(gray_img[1566]), .B2(
        n22694), .O(n21240) );
  OA112S U26746 ( .C1(n29514), .C2(n22251), .A1(n21241), .B1(n21240), .O(
        n21273) );
  INV1S U26747 ( .I(n22853), .O(n22931) );
  ND2S U26748 ( .I1(n22931), .I2(gray_img[1934]), .O(n21252) );
  AOI22S U26749 ( .A1(n22762), .A2(gray_img[398]), .B1(gray_img[1054]), .B2(
        n22935), .O(n21245) );
  AOI22S U26750 ( .A1(n22787), .A2(gray_img[1822]), .B1(gray_img[1286]), .B2(
        n22934), .O(n21244) );
  AOI22S U26751 ( .A1(n22625), .A2(gray_img[262]), .B1(gray_img[782]), .B2(
        n22932), .O(n21243) );
  INV1S U26752 ( .I(gray_img[1798]), .O(n29397) );
  INV1S U26753 ( .I(n22937), .O(n22175) );
  INV1S U26754 ( .I(n22175), .O(n22727) );
  MOAI1S U26755 ( .A1(n22364), .A2(n29397), .B1(n22727), .B2(gray_img[1806]), 
        .O(n21242) );
  AN4B1S U26756 ( .I1(n21245), .I2(n21244), .I3(n21243), .B1(n21242), .O(
        n21251) );
  AOI22S U26757 ( .A1(n15905), .A2(gray_img[278]), .B1(gray_img[1046]), .B2(
        n22929), .O(n21250) );
  ND2S U26758 ( .I1(n15918), .I2(gray_img[150]), .O(n21248) );
  AOI22S U26759 ( .A1(n22735), .A2(gray_img[286]), .B1(gray_img[1542]), .B2(
        n21097), .O(n21247) );
  AOI22S U26760 ( .A1(n22770), .A2(gray_img[1670]), .B1(gray_img[774]), .B2(
        n22513), .O(n21246) );
  ND3S U26761 ( .I1(n21248), .I2(n21247), .I3(n21246), .O(n21249) );
  AN4B1S U26762 ( .I1(n21252), .I2(n21251), .I3(n21250), .B1(n21249), .O(
        n21272) );
  AOI22S U26763 ( .A1(n22888), .A2(gray_img[654]), .B1(gray_img[526]), .B2(
        n22887), .O(n21256) );
  ND2S U26764 ( .I1(n22863), .I2(gray_img[1814]), .O(n21255) );
  AOI22S U26765 ( .A1(n22910), .A2(gray_img[910]), .B1(gray_img[1694]), .B2(
        n22505), .O(n21254) );
  NR2 U26766 ( .I1(n29757), .I2(n22797), .O(n21253) );
  AN4B1S U26767 ( .I1(n21256), .I2(n21255), .I3(n21254), .B1(n21253), .O(
        n21266) );
  AOI22S U26768 ( .A1(n22664), .A2(gray_img[1430]), .B1(gray_img[1174]), .B2(
        n15921), .O(n21265) );
  AOI22S U26769 ( .A1(n22810), .A2(gray_img[646]), .B1(gray_img[390]), .B2(
        n22686), .O(n21264) );
  INV1S U26770 ( .I(gray_img[14]), .O(n23428) );
  ND2S U26771 ( .I1(n22819), .I2(gray_img[926]), .O(n21262) );
  ND2S U26772 ( .I1(n22812), .I2(gray_img[1926]), .O(n21260) );
  AOI22S U26773 ( .A1(gray_img[1182]), .A2(n21090), .B1(gray_img[22]), .B2(
        n22901), .O(n21259) );
  ND2S U26774 ( .I1(gray_img[790]), .I2(n22930), .O(n21258) );
  INV1S U26775 ( .I(gray_img[1310]), .O(n29770) );
  INV1S U26776 ( .I(n21120), .O(n22103) );
  MOAI1S U26777 ( .A1(n29770), .A2(n22103), .B1(gray_img[1942]), .B2(n22679), 
        .O(n21257) );
  AN4B1S U26778 ( .I1(n21260), .I2(n21259), .I3(n21258), .B1(n21257), .O(
        n21261) );
  OAI112HS U26779 ( .C1(n22811), .C2(n23428), .A1(n21262), .B1(n21261), .O(
        n21263) );
  AN4B1S U26780 ( .I1(n21266), .I2(n21265), .I3(n21264), .B1(n21263), .O(
        n21271) );
  ND2S U26781 ( .I1(n22893), .I2(gray_img[6]), .O(n21269) );
  AOI22S U26782 ( .A1(n22828), .A2(gray_img[918]), .B1(gray_img[1558]), .B2(
        n15919), .O(n21268) );
  ND2S U26783 ( .I1(n21137), .I2(gray_img[30]), .O(n21267) );
  ND3S U26784 ( .I1(n21269), .I2(n21268), .I3(n21267), .O(n21270) );
  AN4B1S U26785 ( .I1(n21273), .I2(n21272), .I3(n21271), .B1(n21270), .O(
        n21274) );
  ND3S U26786 ( .I1(n21276), .I2(n21275), .I3(n21274), .O(n21334) );
  NR2 U26787 ( .I1(n30305), .I2(n30307), .O(n22959) );
  INV1S U26788 ( .I(gray_img[366]), .O(n27461) );
  MOAI1S U26789 ( .A1(n22865), .A2(n27461), .B1(n22724), .B2(gray_img[878]), 
        .O(n21281) );
  INV1S U26790 ( .I(gray_img[1134]), .O(n28053) );
  MOAI1S U26791 ( .A1(n22848), .A2(n28053), .B1(n22934), .B2(gray_img[1382]), 
        .O(n21280) );
  INV1S U26792 ( .I(gray_img[1398]), .O(n27915) );
  AOI22S U26793 ( .A1(gray_img[1534]), .A2(n21096), .B1(n21097), .B2(
        gray_img[1638]), .O(n21278) );
  ND2S U26794 ( .I1(n21120), .I2(gray_img[1406]), .O(n21277) );
  OAI112HS U26795 ( .C1(n22797), .C2(n27915), .A1(n21278), .B1(n21277), .O(
        n21279) );
  NR3 U26796 ( .I1(n21281), .I2(n21280), .I3(n21279), .O(n21332) );
  ND2S U26797 ( .I1(n22929), .I2(gray_img[1142]), .O(n21287) );
  AOI22S U26798 ( .A1(n15921), .A2(gray_img[1270]), .B1(gray_img[1654]), .B2(
        n15919), .O(n21286) );
  ND2S U26799 ( .I1(n21152), .I2(gray_img[638]), .O(n21285) );
  AOI22S U26800 ( .A1(n22727), .A2(gray_img[1902]), .B1(gray_img[1774]), .B2(
        n22921), .O(n21283) );
  AOI22S U26801 ( .A1(gray_img[1278]), .A2(n21090), .B1(n22810), .B2(
        gray_img[742]), .O(n21282) );
  ND2S U26802 ( .I1(n21283), .I2(n21282), .O(n21284) );
  AN4B1S U26803 ( .I1(n21287), .I2(n21286), .I3(n21285), .B1(n21284), .O(
        n21331) );
  INV1S U26804 ( .I(gray_img[766]), .O(n26342) );
  MOAI1S U26805 ( .A1(n22803), .A2(n26342), .B1(n22505), .B2(gray_img[1790]), 
        .O(n21290) );
  INV1S U26806 ( .I(gray_img[510]), .O(n27620) );
  MOAI1S U26807 ( .A1(n21288), .A2(n27620), .B1(n22785), .B2(gray_img[382]), 
        .O(n21289) );
  NR2 U26808 ( .I1(n21290), .I2(n21289), .O(n21293) );
  AOI22S U26809 ( .A1(n22888), .A2(gray_img[750]), .B1(gray_img[622]), .B2(
        n22887), .O(n21292) );
  ND2S U26810 ( .I1(n22863), .I2(gray_img[1910]), .O(n21291) );
  ND3S U26811 ( .I1(n21293), .I2(n21292), .I3(n21291), .O(n21309) );
  ND2S U26812 ( .I1(n22893), .I2(gray_img[102]), .O(n21296) );
  BUF1 U26813 ( .I(n22828), .O(n22894) );
  AOI22S U26814 ( .A1(n22619), .A2(gray_img[502]), .B1(gray_img[1014]), .B2(
        n22894), .O(n21295) );
  AOI22S U26815 ( .A1(n22920), .A2(gray_img[758]), .B1(gray_img[1526]), .B2(
        n22664), .O(n21294) );
  ND3S U26816 ( .I1(n21296), .I2(n21295), .I3(n21294), .O(n21308) );
  ND2S U26817 ( .I1(n22896), .I2(gray_img[1782]), .O(n21303) );
  ND2S U26818 ( .I1(n22819), .I2(gray_img[1022]), .O(n21302) );
  ND2S U26819 ( .I1(n22812), .I2(gray_img[2022]), .O(n21301) );
  INV1S U26820 ( .I(n22811), .O(n22900) );
  ND2S U26821 ( .I1(n22900), .I2(gray_img[110]), .O(n21299) );
  AOI22S U26822 ( .A1(gray_img[2038]), .A2(n22679), .B1(gray_img[374]), .B2(
        n15905), .O(n21298) );
  ND2S U26823 ( .I1(gray_img[118]), .I2(n22901), .O(n21297) );
  ND3S U26824 ( .I1(n21299), .I2(n21298), .I3(n21297), .O(n21300) );
  AN4B1S U26825 ( .I1(n21303), .I2(n21302), .I3(n21301), .B1(n21300), .O(
        n21306) );
  AOI22S U26826 ( .A1(n22630), .A2(gray_img[614]), .B1(gray_img[486]), .B2(
        n22686), .O(n21305) );
  AOI22S U26827 ( .A1(n22911), .A2(gray_img[998]), .B1(gray_img[1006]), .B2(
        n22910), .O(n21304) );
  ND3S U26828 ( .I1(n21306), .I2(n21305), .I3(n21304), .O(n21307) );
  NR3 U26829 ( .I1(n21309), .I2(n21308), .I3(n21307), .O(n21316) );
  INV1S U26830 ( .I(n22694), .O(n22618) );
  INV1S U26831 ( .I(n22618), .O(n22918) );
  AOI22S U26832 ( .A1(n22918), .A2(gray_img[1662]), .B1(n21137), .B2(
        gray_img[126]), .O(n21315) );
  ND2S U26833 ( .I1(n22919), .I2(gray_img[2046]), .O(n21314) );
  AOI22S U26834 ( .A1(n22867), .A2(gray_img[894]), .B1(gray_img[254]), .B2(
        n21089), .O(n21312) );
  AOI22S U26835 ( .A1(n22861), .A2(gray_img[1390]), .B1(gray_img[1262]), .B2(
        n22936), .O(n21311) );
  AOI22S U26836 ( .A1(n22656), .A2(gray_img[1646]), .B1(gray_img[1518]), .B2(
        n22369), .O(n21310) );
  ND3S U26837 ( .I1(n21312), .I2(n21311), .I3(n21310), .O(n21313) );
  AN4B1S U26838 ( .I1(n21316), .I2(n21315), .I3(n21314), .B1(n21313), .O(
        n21329) );
  AOI22S U26839 ( .A1(n15915), .A2(gray_img[630]), .B1(gray_img[886]), .B2(
        n22930), .O(n21328) );
  ND2S U26840 ( .I1(n22931), .I2(gray_img[2030]), .O(n21322) );
  AOI22S U26841 ( .A1(n22625), .A2(gray_img[358]), .B1(gray_img[870]), .B2(
        n22513), .O(n21321) );
  AOI22S U26842 ( .A1(n22836), .A2(gray_img[238]), .B1(gray_img[494]), .B2(
        n22862), .O(n21320) );
  AOI22S U26843 ( .A1(n22938), .A2(gray_img[1894]), .B1(gray_img[1126]), .B2(
        n22703), .O(n21318) );
  AOI22S U26844 ( .A1(n22935), .A2(gray_img[1150]), .B1(gray_img[1918]), .B2(
        n22864), .O(n21317) );
  ND2S U26845 ( .I1(n21318), .I2(n21317), .O(n21319) );
  AN4B1S U26846 ( .I1(n21322), .I2(n21321), .I3(n21320), .B1(n21319), .O(
        n21327) );
  ND2S U26847 ( .I1(n15918), .I2(gray_img[246]), .O(n21325) );
  AOI22S U26848 ( .A1(n22770), .A2(gray_img[1766]), .B1(gray_img[1254]), .B2(
        n22838), .O(n21324) );
  AOI22S U26849 ( .A1(n21106), .A2(gray_img[1510]), .B1(gray_img[230]), .B2(
        n22610), .O(n21323) );
  ND3S U26850 ( .I1(n21325), .I2(n21324), .I3(n21323), .O(n21326) );
  AN4B1S U26851 ( .I1(n21329), .I2(n21328), .I3(n21327), .B1(n21326), .O(
        n21330) );
  ND3S U26852 ( .I1(n21332), .I2(n21331), .I3(n21330), .O(n21333) );
  AOI22S U26853 ( .A1(n22784), .A2(n21334), .B1(n22959), .B2(n21333), .O(
        n21335) );
  ND2S U26854 ( .I1(n15918), .I2(gray_img[243]), .O(n21338) );
  AOI22S U26855 ( .A1(n22724), .A2(gray_img[875]), .B1(gray_img[1891]), .B2(
        n22794), .O(n21337) );
  OAI112HS U26856 ( .C1(n22725), .C2(n26392), .A1(n21338), .B1(n21337), .O(
        n21342) );
  INV1S U26857 ( .I(n21089), .O(n21828) );
  AOI22S U26858 ( .A1(gray_img[1275]), .A2(n21090), .B1(n22625), .B2(
        gray_img[355]), .O(n21340) );
  ND2S U26859 ( .I1(n22934), .I2(gray_img[1379]), .O(n21339) );
  OAI112HS U26860 ( .C1(n21828), .C2(n27560), .A1(n21340), .B1(n21339), .O(
        n21341) );
  NR2 U26861 ( .I1(n21342), .I2(n21341), .O(n21399) );
  AOI22S U26862 ( .A1(n22862), .A2(gray_img[491]), .B1(gray_img[1147]), .B2(
        n22935), .O(n21348) );
  ND2S U26863 ( .I1(n22694), .I2(gray_img[1659]), .O(n21345) );
  INV1S U26864 ( .I(n22888), .O(n21884) );
  INV1S U26865 ( .I(n21884), .O(n22657) );
  AOI22S U26866 ( .A1(n22819), .A2(gray_img[1019]), .B1(gray_img[747]), .B2(
        n22657), .O(n21344) );
  ND2S U26867 ( .I1(n22894), .I2(gray_img[1011]), .O(n21343) );
  ND3S U26868 ( .I1(n21345), .I2(n21344), .I3(n21343), .O(n21347) );
  INV1S U26869 ( .I(gray_img[1507]), .O(n27990) );
  MOAI1S U26870 ( .A1(n22718), .A2(n27990), .B1(n22610), .B2(gray_img[227]), 
        .O(n21346) );
  AN3B2S U26871 ( .I1(n21348), .B1(n21347), .B2(n21346), .O(n21398) );
  NR2 U26872 ( .I1(n25852), .I2(n22853), .O(n21353) );
  ND2S U26873 ( .I1(n22929), .I2(gray_img[1139]), .O(n21351) );
  BUF1 U26874 ( .I(n22836), .O(n22933) );
  AOI22S U26875 ( .A1(n22933), .A2(gray_img[235]), .B1(gray_img[1915]), .B2(
        n22787), .O(n21350) );
  AOI22S U26876 ( .A1(n22703), .A2(gray_img[1123]), .B1(gray_img[1259]), .B2(
        n22936), .O(n21349) );
  ND3S U26877 ( .I1(n21351), .I2(n21350), .I3(n21349), .O(n21352) );
  NR2 U26878 ( .I1(n21353), .I2(n21352), .O(n21359) );
  AOI22S U26879 ( .A1(n15905), .A2(gray_img[371]), .B1(gray_img[627]), .B2(
        n15915), .O(n21358) );
  ND2S U26880 ( .I1(n22930), .I2(gray_img[883]), .O(n21356) );
  AOI22S U26881 ( .A1(n21097), .A2(gray_img[1635]), .B1(gray_img[1251]), .B2(
        n22838), .O(n21355) );
  AOI22S U26882 ( .A1(n22513), .A2(gray_img[867]), .B1(gray_img[363]), .B2(
        n22837), .O(n21354) );
  AN3S U26883 ( .I1(n21356), .I2(n21355), .I3(n21354), .O(n21357) );
  ND3S U26884 ( .I1(n21359), .I2(n21358), .I3(n21357), .O(n21396) );
  INV1S U26885 ( .I(gray_img[1771]), .O(n21360) );
  MOAI1S U26886 ( .A1(n22487), .A2(n21360), .B1(n22727), .B2(gray_img[1899]), 
        .O(n21362) );
  INV1S U26887 ( .I(gray_img[1131]), .O(n28047) );
  MOAI1S U26888 ( .A1(n22848), .A2(n28047), .B1(n22861), .B2(gray_img[1387]), 
        .O(n21361) );
  NR2 U26889 ( .I1(n21362), .I2(n21361), .O(n21365) );
  INV1S U26890 ( .I(n22656), .O(n22218) );
  INV1S U26891 ( .I(n22218), .O(n22874) );
  AOI22S U26892 ( .A1(n22874), .A2(gray_img[1643]), .B1(gray_img[1515]), .B2(
        n22369), .O(n21364) );
  ND2S U26893 ( .I1(n21152), .I2(gray_img[635]), .O(n21363) );
  ND3S U26894 ( .I1(n21365), .I2(n21364), .I3(n21363), .O(n21370) );
  ND2S U26895 ( .I1(n22755), .I2(gray_img[2043]), .O(n21368) );
  AOI22S U26896 ( .A1(n22619), .A2(gray_img[499]), .B1(gray_img[755]), .B2(
        n22920), .O(n21367) );
  ND2S U26897 ( .I1(n21137), .I2(gray_img[123]), .O(n21366) );
  ND3S U26898 ( .I1(n21368), .I2(n21367), .I3(n21366), .O(n21369) );
  NR2 U26899 ( .I1(n21370), .I2(n21369), .O(n21394) );
  INV1S U26900 ( .I(gray_img[995]), .O(n26247) );
  AOI22S U26901 ( .A1(n22630), .A2(gray_img[611]), .B1(gray_img[739]), .B2(
        n22909), .O(n21378) );
  INV1S U26902 ( .I(gray_img[107]), .O(n21371) );
  NR2 U26903 ( .I1(n21371), .I2(n22811), .O(n21376) );
  ND2S U26904 ( .I1(n22812), .I2(gray_img[2019]), .O(n21374) );
  AOI22S U26905 ( .A1(gray_img[1531]), .A2(n21096), .B1(gray_img[2035]), .B2(
        n22679), .O(n21373) );
  AOI22S U26906 ( .A1(gray_img[115]), .A2(n22901), .B1(gray_img[1403]), .B2(
        n21120), .O(n21372) );
  ND3S U26907 ( .I1(n21374), .I2(n21373), .I3(n21372), .O(n21375) );
  NR2 U26908 ( .I1(n21376), .I2(n21375), .O(n21377) );
  OAI112HS U26909 ( .C1(n21841), .C2(n26247), .A1(n21378), .B1(n21377), .O(
        n21388) );
  ND2S U26910 ( .I1(n22863), .I2(gray_img[1907]), .O(n21380) );
  BUF1 U26911 ( .I(n22887), .O(n22795) );
  AOI22S U26912 ( .A1(n22686), .A2(gray_img[483]), .B1(gray_img[619]), .B2(
        n22795), .O(n21379) );
  ND2S U26913 ( .I1(n21380), .I2(n21379), .O(n21387) );
  INV1S U26914 ( .I(gray_img[1787]), .O(n25987) );
  MOAI1S U26915 ( .A1(n22882), .A2(n25987), .B1(n22802), .B2(gray_img[1003]), 
        .O(n21382) );
  INV1S U26916 ( .I(gray_img[1395]), .O(n27909) );
  NR2 U26917 ( .I1(n27909), .I2(n22797), .O(n21381) );
  NR2 U26918 ( .I1(n21382), .I2(n21381), .O(n21385) );
  AOI22S U26919 ( .A1(n22883), .A2(gray_img[763]), .B1(gray_img[507]), .B2(
        n22736), .O(n21384) );
  AOI22S U26920 ( .A1(n22735), .A2(gray_img[379]), .B1(gray_img[1763]), .B2(
        n22770), .O(n21383) );
  ND3S U26921 ( .I1(n21385), .I2(n21384), .I3(n21383), .O(n21386) );
  NR3 U26922 ( .I1(n21388), .I2(n21387), .I3(n21386), .O(n21393) );
  ND2S U26923 ( .I1(n22893), .I2(gray_img[99]), .O(n21391) );
  AOI22S U26924 ( .A1(n22796), .A2(gray_img[1779]), .B1(gray_img[1523]), .B2(
        n22664), .O(n21390) );
  AOI22S U26925 ( .A1(n15921), .A2(gray_img[1267]), .B1(gray_img[1651]), .B2(
        n15919), .O(n21389) );
  AN3S U26926 ( .I1(n21391), .I2(n21390), .I3(n21389), .O(n21392) );
  ND3S U26927 ( .I1(n21394), .I2(n21393), .I3(n21392), .O(n21395) );
  NR2 U26928 ( .I1(n21396), .I2(n21395), .O(n21397) );
  AOI22S U26929 ( .A1(n22874), .A2(gray_img[1579]), .B1(n22664), .B2(
        gray_img[1459]), .O(n21403) );
  AOI22S U26930 ( .A1(gray_img[1211]), .A2(n21090), .B1(n22630), .B2(
        gray_img[547]), .O(n21402) );
  AOI22S U26931 ( .A1(n22657), .A2(gray_img[683]), .B1(gray_img[555]), .B2(
        n22887), .O(n21401) );
  INV1S U26932 ( .I(gray_img[1451]), .O(n28966) );
  MOAI1S U26933 ( .A1(n22875), .A2(n28966), .B1(n22881), .B2(gray_img[443]), 
        .O(n21400) );
  AN4B1S U26934 ( .I1(n21403), .I2(n21402), .I3(n21401), .B1(n21400), .O(
        n21449) );
  AOI22S U26935 ( .A1(n22727), .A2(gray_img[1835]), .B1(n22827), .B2(
        gray_img[1587]), .O(n21407) );
  AOI22S U26936 ( .A1(n22762), .A2(gray_img[427]), .B1(n21155), .B2(
        gray_img[1067]), .O(n21406) );
  AOI22S U26937 ( .A1(n22873), .A2(gray_img[955]), .B1(n22610), .B2(
        gray_img[163]), .O(n21405) );
  MOAI1S U26938 ( .A1(n22865), .A2(n27279), .B1(n22724), .B2(gray_img[811]), 
        .O(n21404) );
  AN4B1S U26939 ( .I1(n21407), .I2(n21406), .I3(n21405), .B1(n21404), .O(
        n21448) );
  MOAI1S U26940 ( .A1(n22924), .A2(n27713), .B1(gray_img[1467]), .B2(n21096), 
        .O(n21413) );
  INV1S U26941 ( .I(gray_img[1979]), .O(n23130) );
  NR2 U26942 ( .I1(n23130), .I2(n22251), .O(n21412) );
  ND2S U26943 ( .I1(n22893), .I2(gray_img[35]), .O(n21410) );
  AOI22S U26944 ( .A1(n22936), .A2(gray_img[1195]), .B1(n22894), .B2(
        gray_img[947]), .O(n21409) );
  AOI22S U26945 ( .A1(n22619), .A2(gray_img[435]), .B1(gray_img[691]), .B2(
        n22920), .O(n21408) );
  ND3S U26946 ( .I1(n21410), .I2(n21409), .I3(n21408), .O(n21411) );
  NR3 U26947 ( .I1(n21413), .I2(n21412), .I3(n21411), .O(n21433) );
  INV1S U26948 ( .I(gray_img[1715]), .O(n29213) );
  MOAI1S U26949 ( .A1(n22540), .A2(n29213), .B1(n15921), .B2(gray_img[1203]), 
        .O(n21426) );
  AOI22S U26950 ( .A1(n22566), .A2(gray_img[931]), .B1(gray_img[675]), .B2(
        n22810), .O(n21420) );
  ND2S U26951 ( .I1(n22900), .I2(gray_img[43]), .O(n21417) );
  AOI22S U26952 ( .A1(gray_img[51]), .A2(n22901), .B1(gray_img[1339]), .B2(
        n21120), .O(n21416) );
  ND2S U26953 ( .I1(n22812), .I2(gray_img[1955]), .O(n21415) );
  MOAI1S U26954 ( .A1(n28147), .A2(n22750), .B1(gray_img[1971]), .B2(n22679), 
        .O(n21414) );
  AN4B1S U26955 ( .I1(n21417), .I2(n21416), .I3(n21415), .B1(n21414), .O(
        n21419) );
  ND2S U26956 ( .I1(n22686), .I2(gray_img[419]), .O(n21418) );
  ND3S U26957 ( .I1(n21420), .I2(n21419), .I3(n21418), .O(n21425) );
  AOI22S U26958 ( .A1(n22863), .A2(gray_img[1843]), .B1(gray_img[1331]), .B2(
        n22889), .O(n21423) );
  AOI22S U26959 ( .A1(n22802), .A2(gray_img[939]), .B1(gray_img[1723]), .B2(
        n22505), .O(n21422) );
  AOI22S U26960 ( .A1(n22883), .A2(gray_img[699]), .B1(gray_img[315]), .B2(
        n22735), .O(n21421) );
  ND3S U26961 ( .I1(n21423), .I2(n21422), .I3(n21421), .O(n21424) );
  NR3 U26962 ( .I1(n21426), .I2(n21425), .I3(n21424), .O(n21432) );
  AOI22S U26963 ( .A1(n15905), .A2(gray_img[307]), .B1(gray_img[819]), .B2(
        n22930), .O(n21431) );
  ND2S U26964 ( .I1(n15918), .I2(gray_img[179]), .O(n21429) );
  AOI22S U26965 ( .A1(n22770), .A2(gray_img[1699]), .B1(gray_img[1571]), .B2(
        n21097), .O(n21428) );
  AOI22S U26966 ( .A1(n21106), .A2(gray_img[1443]), .B1(gray_img[1187]), .B2(
        n22838), .O(n21427) );
  ND3S U26967 ( .I1(n21429), .I2(n21428), .I3(n21427), .O(n21430) );
  AN4B1S U26968 ( .I1(n21433), .I2(n21432), .I3(n21431), .B1(n21430), .O(
        n21446) );
  AOI22S U26969 ( .A1(n15915), .A2(gray_img[563]), .B1(gray_img[1075]), .B2(
        n22929), .O(n21439) );
  AOI22S U26970 ( .A1(n22625), .A2(gray_img[291]), .B1(gray_img[803]), .B2(
        n22513), .O(n21438) );
  AOI22S U26971 ( .A1(n22933), .A2(gray_img[171]), .B1(gray_img[1851]), .B2(
        n22864), .O(n21437) );
  AOI22S U26972 ( .A1(n22938), .A2(gray_img[1827]), .B1(gray_img[1315]), .B2(
        n22934), .O(n21435) );
  AOI22S U26973 ( .A1(n22935), .A2(gray_img[1083]), .B1(gray_img[1059]), .B2(
        n22703), .O(n21434) );
  ND2S U26974 ( .I1(n21435), .I2(n21434), .O(n21436) );
  AN4B1S U26975 ( .I1(n21439), .I2(n21438), .I3(n21437), .B1(n21436), .O(
        n21445) );
  ND2S U26976 ( .I1(n22931), .I2(gray_img[1963]), .O(n21444) );
  AOI22S U26977 ( .A1(n21089), .A2(gray_img[187]), .B1(gray_img[1595]), .B2(
        n22918), .O(n21442) );
  AOI22S U26978 ( .A1(n22846), .A2(gray_img[1323]), .B1(gray_img[1707]), .B2(
        n22921), .O(n21441) );
  ND2S U26979 ( .I1(n22867), .I2(gray_img[827]), .O(n21440) );
  ND3S U26980 ( .I1(n21442), .I2(n21441), .I3(n21440), .O(n21443) );
  AN4B1S U26981 ( .I1(n21446), .I2(n21445), .I3(n21444), .B1(n21443), .O(
        n21447) );
  AOI22S U26982 ( .A1(n22959), .A2(n21451), .B1(n22957), .B2(n21450), .O(
        n21560) );
  INV1S U26983 ( .I(gray_img[1691]), .O(n26534) );
  MOAI1S U26984 ( .A1(n22882), .A2(n26534), .B1(n22883), .B2(gray_img[667]), 
        .O(n21457) );
  NR2 U26985 ( .I1(n29751), .I2(n22797), .O(n21456) );
  AOI22S U26986 ( .A1(n22727), .A2(gray_img[1803]), .B1(n22695), .B2(
        gray_img[659]), .O(n21454) );
  AOI22S U26987 ( .A1(gray_img[531]), .A2(n15915), .B1(n22911), .B2(
        gray_img[899]), .O(n21453) );
  ND2S U26988 ( .I1(n22828), .I2(gray_img[915]), .O(n21452) );
  ND3S U26989 ( .I1(n21454), .I2(n21453), .I3(n21452), .O(n21455) );
  NR3 U26990 ( .I1(n21457), .I2(n21456), .I3(n21455), .O(n21503) );
  AOI22S U26991 ( .A1(n22610), .A2(gray_img[131]), .B1(gray_img[1795]), .B2(
        n22794), .O(n21461) );
  AOI22S U26992 ( .A1(n22630), .A2(gray_img[515]), .B1(gray_img[651]), .B2(
        n22657), .O(n21460) );
  AOI22S U26993 ( .A1(gray_img[1563]), .A2(n22694), .B1(n22873), .B2(
        gray_img[923]), .O(n21459) );
  INV1S U26994 ( .I(gray_img[403]), .O(n28738) );
  MOAI1S U26995 ( .A1(n22658), .A2(n28738), .B1(gray_img[1419]), .B2(n22847), 
        .O(n21458) );
  AN4B1S U26996 ( .I1(n21461), .I2(n21460), .I3(n21459), .B1(n21458), .O(
        n21502) );
  INV1S U26997 ( .I(gray_img[1931]), .O(n29404) );
  ND2S U26998 ( .I1(n22929), .I2(gray_img[1043]), .O(n21468) );
  AOI22S U26999 ( .A1(n22837), .A2(gray_img[267]), .B1(gray_img[779]), .B2(
        n22724), .O(n21467) );
  AOI22S U27000 ( .A1(n22933), .A2(gray_img[139]), .B1(gray_img[1051]), .B2(
        n22935), .O(n21466) );
  ND2S U27001 ( .I1(n22930), .I2(gray_img[787]), .O(n21464) );
  AOI22S U27002 ( .A1(n21106), .A2(gray_img[1411]), .B1(gray_img[259]), .B2(
        n22625), .O(n21463) );
  AOI22S U27003 ( .A1(n22513), .A2(gray_img[771]), .B1(gray_img[395]), .B2(
        n22862), .O(n21462) );
  ND3S U27004 ( .I1(n21464), .I2(n21463), .I3(n21462), .O(n21465) );
  AN4B1S U27005 ( .I1(n21468), .I2(n21467), .I3(n21466), .B1(n21465), .O(
        n21474) );
  AOI22S U27006 ( .A1(n22874), .A2(gray_img[1547]), .B1(gray_img[1163]), .B2(
        n22936), .O(n21472) );
  AOI22S U27007 ( .A1(n22934), .A2(gray_img[1283]), .B1(gray_img[1675]), .B2(
        n22921), .O(n21471) );
  AOI22S U27008 ( .A1(n22787), .A2(gray_img[1819]), .B1(gray_img[1027]), .B2(
        n22703), .O(n21470) );
  INV1S U27009 ( .I(gray_img[1035]), .O(n26619) );
  MOAI1S U27010 ( .A1(n22848), .A2(n26619), .B1(n22861), .B2(gray_img[1291]), 
        .O(n21469) );
  AN4B1S U27011 ( .I1(n21472), .I2(n21471), .I3(n21470), .B1(n21469), .O(
        n21473) );
  OAI112HS U27012 ( .C1(n29404), .C2(n22853), .A1(n21474), .B1(n21473), .O(
        n21500) );
  INV1S U27013 ( .I(gray_img[1171]), .O(n29803) );
  MOAI1S U27014 ( .A1(n22058), .A2(n29803), .B1(n15919), .B2(gray_img[1555]), 
        .O(n21485) );
  AOI22S U27015 ( .A1(n22686), .A2(gray_img[387]), .B1(gray_img[907]), .B2(
        n22910), .O(n21482) );
  NR2 U27016 ( .I1(n23422), .I2(n22811), .O(n21479) );
  ND2S U27017 ( .I1(n22812), .I2(gray_img[1923]), .O(n21477) );
  AOI22S U27018 ( .A1(gray_img[1939]), .A2(n22679), .B1(gray_img[1307]), .B2(
        n21120), .O(n21476) );
  AOI22S U27019 ( .A1(gray_img[19]), .A2(n22901), .B1(gray_img[155]), .B2(
        n21089), .O(n21475) );
  NR2 U27020 ( .I1(n21479), .I2(n21478), .O(n21481) );
  ND2S U27021 ( .I1(n22909), .I2(gray_img[643]), .O(n21480) );
  INV1S U27022 ( .I(gray_img[3]), .O(n23436) );
  INV1S U27023 ( .I(n22893), .O(n22125) );
  NR2 U27024 ( .I1(n23436), .I2(n22125), .O(n21483) );
  NR3 U27025 ( .I1(n21485), .I2(n21484), .I3(n21483), .O(n21492) );
  AOI22S U27026 ( .A1(n22770), .A2(gray_img[1667]), .B1(gray_img[1155]), .B2(
        n22838), .O(n21489) );
  ND2S U27027 ( .I1(n22863), .I2(gray_img[1811]), .O(n21488) );
  AOI22S U27028 ( .A1(n22795), .A2(gray_img[523]), .B1(gray_img[411]), .B2(
        n22736), .O(n21487) );
  MOAI1S U27029 ( .A1(n22670), .A2(n26592), .B1(n22785), .B2(gray_img[283]), 
        .O(n21486) );
  AN4B1S U27030 ( .I1(n21489), .I2(n21488), .I3(n21487), .B1(n21486), .O(
        n21491) );
  AOI22S U27031 ( .A1(n15918), .A2(gray_img[147]), .B1(gray_img[275]), .B2(
        n15905), .O(n21490) );
  ND3S U27032 ( .I1(n21492), .I2(n21491), .I3(n21490), .O(n21499) );
  INV1S U27033 ( .I(gray_img[1947]), .O(n29508) );
  AOI22S U27034 ( .A1(n22796), .A2(gray_img[1683]), .B1(gray_img[1427]), .B2(
        n22664), .O(n21494) );
  ND2S U27035 ( .I1(n21137), .I2(gray_img[27]), .O(n21493) );
  AOI22S U27036 ( .A1(n21152), .A2(gray_img[539]), .B1(gray_img[795]), .B2(
        n22813), .O(n21496) );
  AOI22S U27037 ( .A1(n21096), .A2(gray_img[1435]), .B1(gray_img[1179]), .B2(
        n21090), .O(n21495) );
  NR3 U27038 ( .I1(n21500), .I2(n21499), .I3(n21498), .O(n21501) );
  ND3S U27039 ( .I1(n21503), .I2(n21502), .I3(n21501), .O(n21558) );
  INV1S U27040 ( .I(gray_img[1603]), .O(n25670) );
  MOAI1S U27041 ( .A1(n22670), .A2(n25670), .B1(n22887), .B2(gray_img[587]), 
        .O(n21509) );
  INV1S U27042 ( .I(gray_img[1883]), .O(n23251) );
  MOAI1S U27043 ( .A1(n21504), .A2(n23251), .B1(n22625), .B2(gray_img[323]), 
        .O(n21508) );
  INV1S U27044 ( .I(gray_img[603]), .O(n27029) );
  AOI22S U27045 ( .A1(n22630), .A2(gray_img[579]), .B1(gray_img[971]), .B2(
        n22910), .O(n21506) );
  ND2S U27046 ( .I1(n22936), .I2(gray_img[1227]), .O(n21505) );
  OAI112HS U27047 ( .C1(n22750), .C2(n27029), .A1(n21506), .B1(n21505), .O(
        n21507) );
  NR3 U27048 ( .I1(n21509), .I2(n21508), .I3(n21507), .O(n21556) );
  AOI22S U27049 ( .A1(n22895), .A2(gray_img[467]), .B1(gray_img[979]), .B2(
        n22894), .O(n21513) );
  AOI22S U27050 ( .A1(gray_img[1371]), .A2(n21120), .B1(n22881), .B2(
        gray_img[475]), .O(n21512) );
  AOI22S U27051 ( .A1(n22770), .A2(gray_img[1731]), .B1(n22861), .B2(
        gray_img[1355]), .O(n21511) );
  INV1S U27052 ( .I(gray_img[1363]), .O(n28376) );
  MOAI1S U27053 ( .A1(n22797), .A2(n28376), .B1(n15921), .B2(gray_img[1235]), 
        .O(n21510) );
  AN4B1S U27054 ( .I1(n21513), .I2(n21512), .I3(n21511), .B1(n21510), .O(
        n21555) );
  AOI22S U27055 ( .A1(n15905), .A2(gray_img[339]), .B1(gray_img[851]), .B2(
        n22930), .O(n21519) );
  AOI22S U27056 ( .A1(n22810), .A2(gray_img[707]), .B1(gray_img[715]), .B2(
        n22888), .O(n21518) );
  ND2S U27057 ( .I1(n22863), .I2(gray_img[1875]), .O(n21517) );
  INV1S U27058 ( .I(n22392), .O(n22872) );
  AOI22S U27059 ( .A1(n22735), .A2(gray_img[347]), .B1(gray_img[1219]), .B2(
        n22872), .O(n21515) );
  AOI22S U27060 ( .A1(n22786), .A2(gray_img[1755]), .B1(gray_img[731]), .B2(
        n22883), .O(n21514) );
  ND2S U27061 ( .I1(n21515), .I2(n21514), .O(n21516) );
  AN4B1S U27062 ( .I1(n21519), .I2(n21518), .I3(n21517), .B1(n21516), .O(
        n21531) );
  AOI22S U27063 ( .A1(n22796), .A2(gray_img[1747]), .B1(gray_img[1491]), .B2(
        n22664), .O(n21530) );
  ND2S U27064 ( .I1(n22893), .I2(gray_img[67]), .O(n21529) );
  AOI22S U27065 ( .A1(n22566), .A2(gray_img[963]), .B1(gray_img[451]), .B2(
        n22686), .O(n21527) );
  NR2 U27066 ( .I1(n23593), .I2(n22811), .O(n21524) );
  ND2S U27067 ( .I1(n22812), .I2(gray_img[1987]), .O(n21522) );
  AOI22S U27068 ( .A1(gray_img[2003]), .A2(n22679), .B1(gray_img[211]), .B2(
        n15918), .O(n21521) );
  AOI22S U27069 ( .A1(gray_img[1627]), .A2(n22918), .B1(gray_img[83]), .B2(
        n22901), .O(n21520) );
  ND3S U27070 ( .I1(n21522), .I2(n21521), .I3(n21520), .O(n21523) );
  NR2 U27071 ( .I1(n21524), .I2(n21523), .O(n21526) );
  ND2S U27072 ( .I1(n22819), .I2(gray_img[987]), .O(n21525) );
  ND3S U27073 ( .I1(n21527), .I2(n21526), .I3(n21525), .O(n21528) );
  AN4B1S U27074 ( .I1(n21531), .I2(n21530), .I3(n21529), .B1(n21528), .O(
        n21538) );
  AOI22S U27075 ( .A1(n22813), .A2(gray_img[859]), .B1(gray_img[219]), .B2(
        n21089), .O(n21537) );
  AOI22S U27076 ( .A1(n21096), .A2(gray_img[1499]), .B1(gray_img[1243]), .B2(
        n21090), .O(n21536) );
  ND2S U27077 ( .I1(n22755), .I2(gray_img[2011]), .O(n21533) );
  AOI22S U27078 ( .A1(n22695), .A2(gray_img[723]), .B1(gray_img[1619]), .B2(
        n15919), .O(n21532) );
  OAI112HS U27079 ( .C1(n22924), .C2(n21534), .A1(n21533), .B1(n21532), .O(
        n21535) );
  AN4B1S U27080 ( .I1(n21538), .I2(n21537), .I3(n21536), .B1(n21535), .O(
        n21553) );
  ND2S U27081 ( .I1(n22663), .I2(gray_img[1107]), .O(n21545) );
  AOI22S U27082 ( .A1(n22837), .A2(gray_img[331]), .B1(gray_img[843]), .B2(
        n22932), .O(n21544) );
  AOI22S U27083 ( .A1(n22933), .A2(gray_img[203]), .B1(gray_img[1115]), .B2(
        n22935), .O(n21543) );
  ND2S U27084 ( .I1(n15915), .I2(gray_img[595]), .O(n21541) );
  AOI22S U27085 ( .A1(n21106), .A2(gray_img[1475]), .B1(gray_img[195]), .B2(
        n22610), .O(n21540) );
  AOI22S U27086 ( .A1(n22513), .A2(gray_img[835]), .B1(gray_img[459]), .B2(
        n22762), .O(n21539) );
  AN4B1S U27087 ( .I1(n21545), .I2(n21544), .I3(n21543), .B1(n21542), .O(
        n21552) );
  AOI22S U27088 ( .A1(n22794), .A2(gray_img[1859]), .B1(gray_img[1091]), .B2(
        n22703), .O(n21549) );
  AOI22S U27089 ( .A1(n22874), .A2(gray_img[1611]), .B1(gray_img[1867]), .B2(
        n22937), .O(n21548) );
  AOI22S U27090 ( .A1(n22934), .A2(gray_img[1347]), .B1(gray_img[1099]), .B2(
        n21155), .O(n21547) );
  INV1S U27091 ( .I(gray_img[1483]), .O(n23518) );
  MOAI1S U27092 ( .A1(n22875), .A2(n23518), .B1(n22921), .B2(gray_img[1739]), 
        .O(n21546) );
  AN4B1S U27093 ( .I1(n21549), .I2(n21548), .I3(n21547), .B1(n21546), .O(
        n21551) );
  NR2 U27094 ( .I1(n23565), .I2(n22853), .O(n21550) );
  AN4B1S U27095 ( .I1(n21553), .I2(n21552), .I3(n21551), .B1(n21550), .O(
        n21554) );
  ND3S U27096 ( .I1(n21556), .I2(n21555), .I3(n21554), .O(n21557) );
  AOI22S U27097 ( .A1(n22784), .A2(n21558), .B1(n22782), .B2(n21557), .O(
        n21559) );
  ND2S U27098 ( .I1(n15918), .I2(gray_img[244]), .O(n21566) );
  AOI22S U27099 ( .A1(n22864), .A2(gray_img[1916]), .B1(n22695), .B2(
        gray_img[756]), .O(n21565) );
  ND2S U27100 ( .I1(n22863), .I2(gray_img[1908]), .O(n21564) );
  AOI22S U27101 ( .A1(n22566), .A2(gray_img[996]), .B1(gray_img[1004]), .B2(
        n22910), .O(n21562) );
  AOI22S U27102 ( .A1(n22873), .A2(gray_img[1020]), .B1(gray_img[612]), .B2(
        n22630), .O(n21561) );
  ND2S U27103 ( .I1(n21562), .I2(n21561), .O(n21563) );
  AN4B1S U27104 ( .I1(n21566), .I2(n21565), .I3(n21564), .B1(n21563), .O(
        n21612) );
  AOI22S U27105 ( .A1(n22785), .A2(gray_img[380]), .B1(n22938), .B2(
        gray_img[1892]), .O(n21572) );
  ND2S U27106 ( .I1(n22694), .I2(gray_img[1660]), .O(n21569) );
  AOI22S U27107 ( .A1(gray_img[372]), .A2(n15905), .B1(n22657), .B2(
        gray_img[748]), .O(n21568) );
  ND2S U27108 ( .I1(n22727), .I2(gray_img[1900]), .O(n21567) );
  ND3S U27109 ( .I1(n21569), .I2(n21568), .I3(n21567), .O(n21571) );
  INV1S U27110 ( .I(gray_img[1644]), .O(n25786) );
  MOAI1S U27111 ( .A1(n22218), .A2(n25786), .B1(n22847), .B2(gray_img[1516]), 
        .O(n21570) );
  AN3B2S U27112 ( .I1(n21572), .B1(n21571), .B2(n21570), .O(n21611) );
  AOI22S U27113 ( .A1(n21152), .A2(gray_img[636]), .B1(gray_img[252]), .B2(
        n21089), .O(n21575) );
  AOI22S U27114 ( .A1(n22703), .A2(gray_img[1124]), .B1(gray_img[1772]), .B2(
        n22921), .O(n21574) );
  AOI22S U27115 ( .A1(n22846), .A2(gray_img[1388]), .B1(gray_img[1260]), .B2(
        n22936), .O(n21573) );
  ND3S U27116 ( .I1(n21575), .I2(n21574), .I3(n21573), .O(n21577) );
  INV1S U27117 ( .I(n21096), .O(n22493) );
  INV1S U27118 ( .I(gray_img[1532]), .O(n27898) );
  MOAI1S U27119 ( .A1(n22493), .A2(n27898), .B1(n21120), .B2(gray_img[1404]), 
        .O(n21576) );
  AO112S U27120 ( .C1(gray_img[2044]), .C2(n22919), .A1(n21577), .B1(n21576), 
        .O(n21609) );
  INV1S U27121 ( .I(gray_img[100]), .O(n27414) );
  AOI22S U27122 ( .A1(n22664), .A2(gray_img[1524]), .B1(gray_img[1652]), .B2(
        n15919), .O(n21581) );
  ND2S U27123 ( .I1(n21137), .I2(gray_img[124]), .O(n21580) );
  AOI22S U27124 ( .A1(n21155), .A2(gray_img[1132]), .B1(n22619), .B2(
        gray_img[500]), .O(n21579) );
  INV1S U27125 ( .I(gray_img[1780]), .O(n26002) );
  MOAI1S U27126 ( .A1(n22540), .A2(n26002), .B1(n22828), .B2(gray_img[1012]), 
        .O(n21578) );
  AN4B1S U27127 ( .I1(n21581), .I2(n21580), .I3(n21579), .B1(n21578), .O(
        n21594) );
  ND2S U27128 ( .I1(n22889), .I2(gray_img[1396]), .O(n21592) );
  AOI22S U27129 ( .A1(n22686), .A2(gray_img[484]), .B1(gray_img[620]), .B2(
        n22887), .O(n21591) );
  ND2S U27130 ( .I1(n15921), .I2(gray_img[1268]), .O(n21590) );
  ND2S U27131 ( .I1(n22909), .I2(gray_img[740]), .O(n21588) );
  AOI22S U27132 ( .A1(gray_img[1140]), .A2(n22929), .B1(gray_img[892]), .B2(
        n22813), .O(n21585) );
  AOI22S U27133 ( .A1(gray_img[2036]), .A2(n22679), .B1(gray_img[1276]), .B2(
        n21090), .O(n21584) );
  ND2S U27134 ( .I1(gray_img[116]), .I2(n22901), .O(n21583) );
  NR2 U27135 ( .I1(n25842), .I2(n22904), .O(n21582) );
  AN4B1S U27136 ( .I1(n21585), .I2(n21584), .I3(n21583), .B1(n21582), .O(
        n21587) );
  ND2S U27137 ( .I1(n22900), .I2(gray_img[108]), .O(n21586) );
  ND3S U27138 ( .I1(n21588), .I2(n21587), .I3(n21586), .O(n21589) );
  AN4B1S U27139 ( .I1(n21592), .I2(n21591), .I3(n21590), .B1(n21589), .O(
        n21593) );
  OAI112HS U27140 ( .C1(n27414), .C2(n22125), .A1(n21594), .B1(n21593), .O(
        n21608) );
  AOI22S U27141 ( .A1(n22933), .A2(gray_img[236]), .B1(gray_img[492]), .B2(
        n22762), .O(n21598) );
  AOI22S U27142 ( .A1(n22935), .A2(gray_img[1148]), .B1(gray_img[1380]), .B2(
        n22934), .O(n21597) );
  AOI22S U27143 ( .A1(n22513), .A2(gray_img[868]), .B1(gray_img[228]), .B2(
        n22610), .O(n21596) );
  INV1S U27144 ( .I(gray_img[364]), .O(n27457) );
  MOAI1S U27145 ( .A1(n22865), .A2(n27457), .B1(n22932), .B2(gray_img[876]), 
        .O(n21595) );
  AN4B1S U27146 ( .I1(n21598), .I2(n21597), .I3(n21596), .B1(n21595), .O(
        n21599) );
  OA12S U27147 ( .B1(n25854), .B2(n22853), .A1(n21599), .O(n21606) );
  AOI22S U27148 ( .A1(n22736), .A2(gray_img[508]), .B1(gray_img[1636]), .B2(
        n21097), .O(n21603) );
  AOI22S U27149 ( .A1(n22872), .A2(gray_img[1252]), .B1(gray_img[356]), .B2(
        n22625), .O(n21602) );
  AOI22S U27150 ( .A1(n22786), .A2(gray_img[1788]), .B1(gray_img[764]), .B2(
        n22883), .O(n21601) );
  INV1S U27151 ( .I(gray_img[1508]), .O(n27992) );
  MOAI1S U27152 ( .A1(n22718), .A2(n27992), .B1(n22770), .B2(gray_img[1764]), 
        .O(n21600) );
  AN4B1S U27153 ( .I1(n21603), .I2(n21602), .I3(n21601), .B1(n21600), .O(
        n21605) );
  AOI22S U27154 ( .A1(n15915), .A2(gray_img[628]), .B1(gray_img[884]), .B2(
        n22930), .O(n21604) );
  ND3S U27155 ( .I1(n21606), .I2(n21605), .I3(n21604), .O(n21607) );
  NR3 U27156 ( .I1(n21609), .I2(n21608), .I3(n21607), .O(n21610) );
  ND3S U27157 ( .I1(n21612), .I2(n21611), .I3(n21610), .O(n21664) );
  AOI22S U27158 ( .A1(n21155), .A2(gray_img[1100]), .B1(n22863), .B2(
        gray_img[1876]), .O(n21616) );
  AOI22S U27159 ( .A1(n22630), .A2(gray_img[580]), .B1(gray_img[348]), .B2(
        n22785), .O(n21615) );
  AOI22S U27160 ( .A1(n22938), .A2(gray_img[1860]), .B1(gray_img[1092]), .B2(
        n22703), .O(n21614) );
  INV1S U27161 ( .I(gray_img[1604]), .O(n25672) );
  MOAI1S U27162 ( .A1(n22670), .A2(n25672), .B1(n22625), .B2(gray_img[324]), 
        .O(n21613) );
  AN4B1S U27163 ( .I1(n21616), .I2(n21615), .I3(n21614), .B1(n21613), .O(
        n21662) );
  AOI22S U27164 ( .A1(n22846), .A2(gray_img[1356]), .B1(n22920), .B2(
        gray_img[724]), .O(n21620) );
  AOI22S U27165 ( .A1(n22873), .A2(gray_img[988]), .B1(n22770), .B2(
        gray_img[1732]), .O(n21619) );
  AOI22S U27166 ( .A1(n21106), .A2(gray_img[1476]), .B1(gray_img[332]), .B2(
        n22837), .O(n21618) );
  INV1S U27167 ( .I(gray_img[604]), .O(n27031) );
  MOAI1S U27168 ( .A1(n27031), .A2(n22750), .B1(n21096), .B2(gray_img[1500]), 
        .O(n21617) );
  AN4B1S U27169 ( .I1(n21620), .I2(n21619), .I3(n21618), .B1(n21617), .O(
        n21661) );
  AOI22S U27170 ( .A1(n22664), .A2(gray_img[1492]), .B1(gray_img[1620]), .B2(
        n15919), .O(n21630) );
  ND2S U27171 ( .I1(n22810), .I2(gray_img[708]), .O(n21627) );
  ND2S U27172 ( .I1(n22900), .I2(gray_img[76]), .O(n21626) );
  ND2S U27173 ( .I1(n22812), .I2(gray_img[1988]), .O(n21625) );
  AOI22S U27174 ( .A1(gray_img[2004]), .A2(n22679), .B1(gray_img[212]), .B2(
        n15918), .O(n21623) );
  AOI22S U27175 ( .A1(gray_img[1372]), .A2(n21120), .B1(gray_img[596]), .B2(
        n15915), .O(n21622) );
  ND2S U27176 ( .I1(gray_img[84]), .I2(n22901), .O(n21621) );
  ND3S U27177 ( .I1(n21623), .I2(n21622), .I3(n21621), .O(n21624) );
  AN4B1S U27178 ( .I1(n21627), .I2(n21626), .I3(n21625), .B1(n21624), .O(
        n21629) );
  AOI22S U27179 ( .A1(n22566), .A2(gray_img[964]), .B1(gray_img[452]), .B2(
        n22686), .O(n21628) );
  ND3S U27180 ( .I1(n21630), .I2(n21629), .I3(n21628), .O(n21640) );
  ND2S U27181 ( .I1(n22893), .I2(gray_img[68]), .O(n21633) );
  AOI22S U27182 ( .A1(n22895), .A2(gray_img[468]), .B1(gray_img[980]), .B2(
        n22828), .O(n21632) );
  AOI22S U27183 ( .A1(n22896), .A2(gray_img[1748]), .B1(gray_img[1236]), .B2(
        n15921), .O(n21631) );
  ND3S U27184 ( .I1(n21633), .I2(n21632), .I3(n21631), .O(n21639) );
  INV1S U27185 ( .I(gray_img[1364]), .O(n28378) );
  AOI22S U27186 ( .A1(n22888), .A2(gray_img[716]), .B1(gray_img[588]), .B2(
        n22795), .O(n21634) );
  OA12S U27187 ( .B1(n28378), .B2(n22797), .A1(n21634), .O(n21637) );
  AOI22S U27188 ( .A1(n22802), .A2(gray_img[972]), .B1(gray_img[1756]), .B2(
        n22505), .O(n21636) );
  AOI22S U27189 ( .A1(n22883), .A2(gray_img[732]), .B1(gray_img[476]), .B2(
        n22736), .O(n21635) );
  NR3 U27190 ( .I1(n21640), .I2(n21639), .I3(n21638), .O(n21646) );
  AOI22S U27191 ( .A1(n21090), .A2(gray_img[1244]), .B1(n21137), .B2(
        gray_img[92]), .O(n21645) );
  ND2S U27192 ( .I1(n22755), .I2(gray_img[2012]), .O(n21644) );
  INV1S U27193 ( .I(gray_img[860]), .O(n23072) );
  AOI22S U27194 ( .A1(n21089), .A2(gray_img[220]), .B1(gray_img[1628]), .B2(
        n22918), .O(n21642) );
  AOI22S U27195 ( .A1(n22847), .A2(gray_img[1484]), .B1(gray_img[1740]), .B2(
        n22921), .O(n21641) );
  OAI112HS U27196 ( .C1(n22725), .C2(n23072), .A1(n21642), .B1(n21641), .O(
        n21643) );
  AN4B1S U27197 ( .I1(n21646), .I2(n21645), .I3(n21644), .B1(n21643), .O(
        n21659) );
  AOI22S U27198 ( .A1(n15905), .A2(gray_img[340]), .B1(gray_img[852]), .B2(
        n22930), .O(n21658) );
  ND2S U27199 ( .I1(n22931), .I2(gray_img[1996]), .O(n21652) );
  AOI22S U27200 ( .A1(n22933), .A2(gray_img[204]), .B1(gray_img[460]), .B2(
        n22862), .O(n21651) );
  AOI22S U27201 ( .A1(n22935), .A2(gray_img[1116]), .B1(gray_img[1884]), .B2(
        n22864), .O(n21650) );
  AOI22S U27202 ( .A1(n22874), .A2(gray_img[1612]), .B1(gray_img[1228]), .B2(
        n22936), .O(n21648) );
  AOI22S U27203 ( .A1(n22934), .A2(gray_img[1348]), .B1(gray_img[1868]), .B2(
        n22937), .O(n21647) );
  ND2S U27204 ( .I1(n21648), .I2(n21647), .O(n21649) );
  AN4B1S U27205 ( .I1(n21652), .I2(n21651), .I3(n21650), .B1(n21649), .O(
        n21657) );
  ND2S U27206 ( .I1(n22663), .I2(gray_img[1108]), .O(n21655) );
  AOI22S U27207 ( .A1(n22872), .A2(gray_img[1220]), .B1(gray_img[836]), .B2(
        n22513), .O(n21654) );
  AOI22S U27208 ( .A1(n22610), .A2(gray_img[196]), .B1(gray_img[844]), .B2(
        n22932), .O(n21653) );
  ND3S U27209 ( .I1(n21655), .I2(n21654), .I3(n21653), .O(n21656) );
  AN4B1S U27210 ( .I1(n21659), .I2(n21658), .I3(n21657), .B1(n21656), .O(
        n21660) );
  AOI22S U27211 ( .A1(n22959), .A2(n21664), .B1(n22782), .B2(n21663), .O(
        n21775) );
  ND2S U27212 ( .I1(n21090), .I2(gray_img[1180]), .O(n21669) );
  AOI22S U27213 ( .A1(n22932), .A2(gray_img[780]), .B1(n22847), .B2(
        gray_img[1420]), .O(n21668) );
  AOI22S U27214 ( .A1(n22513), .A2(gray_img[772]), .B1(gray_img[132]), .B2(
        n22610), .O(n21667) );
  INV1S U27215 ( .I(gray_img[1300]), .O(n29753) );
  AOI22S U27216 ( .A1(gray_img[788]), .A2(n22930), .B1(n22566), .B2(
        gray_img[900]), .O(n21665) );
  OAI12HS U27217 ( .B1(n22797), .B2(n29753), .A1(n21665), .O(n21666) );
  AN4B1S U27218 ( .I1(n21669), .I2(n21668), .I3(n21667), .B1(n21666), .O(
        n21721) );
  AOI22S U27219 ( .A1(n22934), .A2(gray_img[1284]), .B1(gray_img[1164]), .B2(
        n22936), .O(n21674) );
  INV1S U27220 ( .I(gray_img[1676]), .O(n26581) );
  ND2S U27221 ( .I1(n15905), .I2(gray_img[276]), .O(n21671) );
  AOI22S U27222 ( .A1(n22819), .A2(gray_img[924]), .B1(gray_img[388]), .B2(
        n22686), .O(n21670) );
  OAI112HS U27223 ( .C1(n22487), .C2(n26581), .A1(n21671), .B1(n21670), .O(
        n21673) );
  MOAI1S U27224 ( .A1(n22392), .A2(n26633), .B1(n22836), .B2(gray_img[140]), 
        .O(n21672) );
  AN3B2S U27225 ( .I1(n21674), .B1(n21673), .B2(n21672), .O(n21720) );
  ND2S U27226 ( .I1(n15918), .I2(gray_img[148]), .O(n21677) );
  AOI22S U27227 ( .A1(n21097), .A2(gray_img[1540]), .B1(gray_img[260]), .B2(
        n22625), .O(n21676) );
  AOI22S U27228 ( .A1(n22837), .A2(gray_img[268]), .B1(gray_img[396]), .B2(
        n22862), .O(n21675) );
  ND3S U27229 ( .I1(n21677), .I2(n21676), .I3(n21675), .O(n21687) );
  ND2S U27230 ( .I1(n22929), .I2(gray_img[1044]), .O(n21680) );
  AOI22S U27231 ( .A1(n22935), .A2(gray_img[1052]), .B1(gray_img[1820]), .B2(
        n22787), .O(n21679) );
  AOI22S U27232 ( .A1(n22794), .A2(gray_img[1796]), .B1(gray_img[1028]), .B2(
        n22703), .O(n21678) );
  ND3S U27233 ( .I1(n21680), .I2(n21679), .I3(n21678), .O(n21686) );
  INV1S U27234 ( .I(gray_img[1292]), .O(n29662) );
  MOAI1S U27235 ( .A1(n22031), .A2(n29662), .B1(n22656), .B2(gray_img[1548]), 
        .O(n21682) );
  INV1S U27236 ( .I(gray_img[1036]), .O(n26621) );
  MOAI1S U27237 ( .A1(n22848), .A2(n26621), .B1(n22727), .B2(gray_img[1804]), 
        .O(n21681) );
  NR2 U27238 ( .I1(n21682), .I2(n21681), .O(n21684) );
  AOI22S U27239 ( .A1(n21152), .A2(gray_img[540]), .B1(gray_img[796]), .B2(
        n22813), .O(n21683) );
  OAI112HS U27240 ( .C1(n22853), .C2(n29406), .A1(n21684), .B1(n21683), .O(
        n21685) );
  NR3 U27241 ( .I1(n21687), .I2(n21686), .I3(n21685), .O(n21718) );
  ND2S U27242 ( .I1(n15919), .I2(gray_img[1556]), .O(n21694) );
  ND2S U27243 ( .I1(n22812), .I2(gray_img[1924]), .O(n21691) );
  AOI22S U27244 ( .A1(gray_img[1940]), .A2(n22679), .B1(gray_img[532]), .B2(
        n15915), .O(n21690) );
  ND2S U27245 ( .I1(gray_img[20]), .I2(n22901), .O(n21689) );
  INV1S U27246 ( .I(gray_img[12]), .O(n23424) );
  NR2 U27247 ( .I1(n23424), .I2(n22811), .O(n21688) );
  AN4B1S U27248 ( .I1(n21691), .I2(n21690), .I3(n21689), .B1(n21688), .O(
        n21693) );
  ND2S U27249 ( .I1(n22909), .I2(gray_img[644]), .O(n21692) );
  AN3S U27250 ( .I1(n21694), .I2(n21693), .I3(n21692), .O(n21697) );
  AOI22S U27251 ( .A1(n22630), .A2(gray_img[516]), .B1(gray_img[908]), .B2(
        n22910), .O(n21696) );
  AOI22S U27252 ( .A1(n22888), .A2(gray_img[652]), .B1(gray_img[524]), .B2(
        n22887), .O(n21695) );
  ND3S U27253 ( .I1(n21697), .I2(n21696), .I3(n21695), .O(n21709) );
  INV1S U27254 ( .I(gray_img[668]), .O(n21698) );
  MOAI1S U27255 ( .A1(n22803), .A2(n21698), .B1(n22785), .B2(gray_img[284]), 
        .O(n21700) );
  INV1S U27256 ( .I(gray_img[1412]), .O(n29650) );
  MOAI1S U27257 ( .A1(n22718), .A2(n29650), .B1(n22770), .B2(gray_img[1668]), 
        .O(n21699) );
  NR2 U27258 ( .I1(n21700), .I2(n21699), .O(n21703) );
  AOI22S U27259 ( .A1(n22786), .A2(gray_img[1692]), .B1(gray_img[412]), .B2(
        n22736), .O(n21702) );
  ND2S U27260 ( .I1(n22863), .I2(gray_img[1812]), .O(n21701) );
  ND3S U27261 ( .I1(n21703), .I2(n21702), .I3(n21701), .O(n21708) );
  ND2S U27262 ( .I1(n22893), .I2(gray_img[4]), .O(n21706) );
  AOI22S U27263 ( .A1(n22695), .A2(gray_img[660]), .B1(gray_img[1684]), .B2(
        n22896), .O(n21705) );
  AOI22S U27264 ( .A1(n22664), .A2(gray_img[1428]), .B1(gray_img[1172]), .B2(
        n15921), .O(n21704) );
  NR3 U27265 ( .I1(n21709), .I2(n21708), .I3(n21707), .O(n21717) );
  INV1S U27266 ( .I(gray_img[156]), .O(n27870) );
  MOAI1S U27267 ( .A1(n27870), .A2(n21828), .B1(n22694), .B2(gray_img[1564]), 
        .O(n21715) );
  INV1S U27268 ( .I(gray_img[1308]), .O(n29766) );
  MOAI1S U27269 ( .A1(n22103), .A2(n29766), .B1(n21096), .B2(gray_img[1436]), 
        .O(n21714) );
  ND2S U27270 ( .I1(n22919), .I2(gray_img[1948]), .O(n21712) );
  AOI22S U27271 ( .A1(n22895), .A2(gray_img[404]), .B1(gray_img[916]), .B2(
        n22894), .O(n21711) );
  ND2S U27272 ( .I1(n21137), .I2(gray_img[28]), .O(n21710) );
  ND3S U27273 ( .I1(n21712), .I2(n21711), .I3(n21710), .O(n21713) );
  NR3 U27274 ( .I1(n21715), .I2(n21714), .I3(n21713), .O(n21716) );
  AN3S U27275 ( .I1(n21718), .I2(n21717), .I3(n21716), .O(n21719) );
  AOI22S U27276 ( .A1(n22727), .A2(gray_img[1836]), .B1(n22664), .B2(
        gray_img[1460]), .O(n21725) );
  AOI22S U27277 ( .A1(gray_img[1212]), .A2(n21090), .B1(n22686), .B2(
        gray_img[420]), .O(n21724) );
  AOI22S U27278 ( .A1(n22883), .A2(gray_img[700]), .B1(gray_img[1572]), .B2(
        n21097), .O(n21723) );
  INV1S U27279 ( .I(gray_img[300]), .O(n27281) );
  MOAI1S U27280 ( .A1(n27281), .A2(n22865), .B1(n22703), .B2(gray_img[1060]), 
        .O(n21722) );
  AN4B1S U27281 ( .I1(n21725), .I2(n21724), .I3(n21723), .B1(n21722), .O(
        n21771) );
  AOI22S U27282 ( .A1(n22934), .A2(gray_img[1316]), .B1(gray_img[1580]), .B2(
        n22656), .O(n21729) );
  AOI22S U27283 ( .A1(n21106), .A2(gray_img[1444]), .B1(gray_img[1852]), .B2(
        n22787), .O(n21728) );
  AOI22S U27284 ( .A1(n22810), .A2(gray_img[676]), .B1(gray_img[444]), .B2(
        n22881), .O(n21727) );
  INV1S U27285 ( .I(gray_img[1708]), .O(n29102) );
  MOAI1S U27286 ( .A1(n29102), .A2(n22487), .B1(n22828), .B2(gray_img[948]), 
        .O(n21726) );
  AN4B1S U27287 ( .I1(n21729), .I2(n21728), .I3(n21727), .B1(n21726), .O(
        n21770) );
  ND2S U27288 ( .I1(n15918), .I2(gray_img[180]), .O(n21732) );
  AOI22S U27289 ( .A1(n22735), .A2(gray_img[316]), .B1(gray_img[1700]), .B2(
        n22770), .O(n21731) );
  AOI22S U27290 ( .A1(n22872), .A2(gray_img[1188]), .B1(gray_img[804]), .B2(
        n22513), .O(n21730) );
  INV1S U27291 ( .I(gray_img[308]), .O(n26507) );
  MOAI1S U27292 ( .A1(n22383), .A2(n26507), .B1(n15915), .B2(gray_img[564]), 
        .O(n21747) );
  ND2S U27293 ( .I1(n22863), .I2(gray_img[1844]), .O(n21736) );
  ND2S U27294 ( .I1(n22889), .I2(gray_img[1332]), .O(n21735) );
  AOI22S U27295 ( .A1(n22802), .A2(gray_img[940]), .B1(gray_img[684]), .B2(
        n22657), .O(n21734) );
  INV1S U27296 ( .I(gray_img[1724]), .O(n29203) );
  MOAI1S U27297 ( .A1(n22882), .A2(n29203), .B1(n22795), .B2(gray_img[556]), 
        .O(n21733) );
  AN4B1S U27298 ( .I1(n21736), .I2(n21735), .I3(n21734), .B1(n21733), .O(
        n21745) );
  AOI22S U27299 ( .A1(n22630), .A2(gray_img[548]), .B1(gray_img[932]), .B2(
        n22566), .O(n21742) );
  ND2S U27300 ( .I1(n22819), .I2(gray_img[956]), .O(n21741) );
  ND2S U27301 ( .I1(n22900), .I2(gray_img[44]), .O(n21740) );
  AOI22S U27302 ( .A1(gray_img[1468]), .A2(n21096), .B1(gray_img[1972]), .B2(
        n22679), .O(n21738) );
  AOI22S U27303 ( .A1(gray_img[52]), .A2(n22901), .B1(gray_img[1596]), .B2(
        n22918), .O(n21737) );
  OAI112HS U27304 ( .C1(n22904), .C2(n26662), .A1(n21738), .B1(n21737), .O(
        n21739) );
  AN4B1S U27305 ( .I1(n21742), .I2(n21741), .I3(n21740), .B1(n21739), .O(
        n21744) );
  AOI22S U27306 ( .A1(n15921), .A2(gray_img[1204]), .B1(gray_img[1588]), .B2(
        n15919), .O(n21743) );
  NR3 U27307 ( .I1(n21748), .I2(n21747), .I3(n21746), .O(n21755) );
  AOI22S U27308 ( .A1(n21120), .A2(gray_img[1340]), .B1(n21137), .B2(
        gray_img[60]), .O(n21754) );
  ND2S U27309 ( .I1(n22919), .I2(gray_img[1980]), .O(n21753) );
  ND2S U27310 ( .I1(n22893), .I2(gray_img[36]), .O(n21751) );
  AOI22S U27311 ( .A1(n22861), .A2(gray_img[1324]), .B1(n22619), .B2(
        gray_img[436]), .O(n21750) );
  AOI22S U27312 ( .A1(n22695), .A2(gray_img[692]), .B1(gray_img[1716]), .B2(
        n22896), .O(n21749) );
  ND3S U27313 ( .I1(n21751), .I2(n21750), .I3(n21749), .O(n21752) );
  AN4B1S U27314 ( .I1(n21755), .I2(n21754), .I3(n21753), .B1(n21752), .O(
        n21768) );
  ND2S U27315 ( .I1(n22663), .I2(gray_img[1076]), .O(n21761) );
  AOI22S U27316 ( .A1(n22724), .A2(gray_img[812]), .B1(gray_img[1084]), .B2(
        n22935), .O(n21760) );
  AOI22S U27317 ( .A1(n22794), .A2(gray_img[1828]), .B1(gray_img[1452]), .B2(
        n22369), .O(n21759) );
  INV1S U27318 ( .I(gray_img[572]), .O(n28149) );
  AOI22S U27319 ( .A1(n22813), .A2(gray_img[828]), .B1(gray_img[188]), .B2(
        n21089), .O(n21757) );
  AOI22S U27320 ( .A1(n21155), .A2(gray_img[1068]), .B1(gray_img[1196]), .B2(
        n22936), .O(n21756) );
  OAI112HS U27321 ( .C1(n22750), .C2(n28149), .A1(n21757), .B1(n21756), .O(
        n21758) );
  AN4B1S U27322 ( .I1(n21761), .I2(n21760), .I3(n21759), .B1(n21758), .O(
        n21767) );
  ND2S U27323 ( .I1(n22931), .I2(gray_img[1964]), .O(n21766) );
  ND2S U27324 ( .I1(n22930), .I2(gray_img[820]), .O(n21764) );
  AOI22S U27325 ( .A1(n22625), .A2(gray_img[292]), .B1(gray_img[164]), .B2(
        n22610), .O(n21763) );
  AOI22S U27326 ( .A1(n22933), .A2(gray_img[172]), .B1(gray_img[428]), .B2(
        n22762), .O(n21762) );
  ND3S U27327 ( .I1(n21764), .I2(n21763), .I3(n21762), .O(n21765) );
  AN4B1S U27328 ( .I1(n21768), .I2(n21767), .I3(n21766), .B1(n21765), .O(
        n21769) );
  AOI22S U27329 ( .A1(n22784), .A2(n21773), .B1(n22957), .B2(n21772), .O(
        n21774) );
  INV1S U27330 ( .I(gray_img[1183]), .O(n29799) );
  INV1S U27331 ( .I(n21090), .O(n22789) );
  NR2 U27332 ( .I1(n29799), .I2(n22789), .O(n21781) );
  INV1S U27333 ( .I(gray_img[1799]), .O(n29399) );
  MOAI1S U27334 ( .A1(n22364), .A2(n29399), .B1(n22864), .B2(gray_img[1823]), 
        .O(n21780) );
  ND2S U27335 ( .I1(n15918), .I2(gray_img[151]), .O(n21778) );
  AOI22S U27336 ( .A1(n22802), .A2(gray_img[911]), .B1(gray_img[1159]), .B2(
        n22838), .O(n21777) );
  AOI22S U27337 ( .A1(n22625), .A2(gray_img[263]), .B1(gray_img[783]), .B2(
        n22932), .O(n21776) );
  ND3S U27338 ( .I1(n21778), .I2(n21777), .I3(n21776), .O(n21779) );
  NR3 U27339 ( .I1(n21781), .I2(n21780), .I3(n21779), .O(n21827) );
  ND2S U27340 ( .I1(n22930), .I2(gray_img[791]), .O(n21786) );
  AOI22S U27341 ( .A1(n22861), .A2(gray_img[1295]), .B1(gray_img[1167]), .B2(
        n22936), .O(n21785) );
  AOI22S U27342 ( .A1(n22770), .A2(gray_img[1671]), .B1(gray_img[143]), .B2(
        n22836), .O(n21784) );
  MOAI1S U27343 ( .A1(n22670), .A2(n26600), .B1(n22505), .B2(gray_img[1695]), 
        .O(n21782) );
  AO12S U27344 ( .B1(gray_img[1431]), .B2(n22664), .A1(n21782), .O(n21783) );
  AN4B1S U27345 ( .I1(n21786), .I2(n21785), .I3(n21784), .B1(n21783), .O(
        n21826) );
  INV1S U27346 ( .I(gray_img[1039]), .O(n26627) );
  MOAI1S U27347 ( .A1(n22848), .A2(n26627), .B1(n22847), .B2(gray_img[1423]), 
        .O(n21789) );
  INV1S U27348 ( .I(gray_img[1679]), .O(n26587) );
  MOAI1S U27349 ( .A1(n22487), .A2(n26587), .B1(n22656), .B2(gray_img[1551]), 
        .O(n21788) );
  INV1S U27350 ( .I(gray_img[543]), .O(n29080) );
  MOAI1S U27351 ( .A1(n22750), .A2(n29080), .B1(n22813), .B2(gray_img[799]), 
        .O(n21787) );
  NR3 U27352 ( .I1(n21789), .I2(n21788), .I3(n21787), .O(n21791) );
  AOI22S U27353 ( .A1(n21096), .A2(gray_img[1439]), .B1(gray_img[1567]), .B2(
        n22694), .O(n21790) );
  OAI112HS U27354 ( .C1(n22251), .C2(n29516), .A1(n21791), .B1(n21790), .O(
        n21824) );
  ND2S U27355 ( .I1(n15905), .I2(gray_img[279]), .O(n21798) );
  AOI22S U27356 ( .A1(n22735), .A2(gray_img[287]), .B1(gray_img[415]), .B2(
        n22736), .O(n21797) );
  AOI22S U27357 ( .A1(n22883), .A2(gray_img[671]), .B1(gray_img[1415]), .B2(
        n21106), .O(n21796) );
  AOI22S U27358 ( .A1(n22863), .A2(gray_img[1815]), .B1(gray_img[1303]), .B2(
        n22889), .O(n21794) );
  AOI22S U27359 ( .A1(n22630), .A2(gray_img[519]), .B1(gray_img[647]), .B2(
        n22909), .O(n21793) );
  AOI22S U27360 ( .A1(n22888), .A2(gray_img[655]), .B1(gray_img[527]), .B2(
        n22887), .O(n21792) );
  AN4B1S U27361 ( .I1(n21798), .I2(n21797), .I3(n21796), .B1(n21795), .O(
        n21806) );
  AOI22S U27362 ( .A1(n22703), .A2(gray_img[1031]), .B1(gray_img[1807]), .B2(
        n22937), .O(n21803) );
  AOI22S U27363 ( .A1(n22935), .A2(gray_img[1055]), .B1(gray_img[1287]), .B2(
        n22934), .O(n21802) );
  AOI22S U27364 ( .A1(n22513), .A2(gray_img[775]), .B1(gray_img[135]), .B2(
        n22610), .O(n21801) );
  MOAI1S U27365 ( .A1(n22865), .A2(n21799), .B1(n22762), .B2(gray_img[399]), 
        .O(n21800) );
  AN4B1S U27366 ( .I1(n21803), .I2(n21802), .I3(n21801), .B1(n21800), .O(
        n21805) );
  ND2S U27367 ( .I1(n22931), .I2(gray_img[1935]), .O(n21804) );
  ND3S U27368 ( .I1(n21806), .I2(n21805), .I3(n21804), .O(n21823) );
  AOI22S U27369 ( .A1(n21120), .A2(gray_img[1311]), .B1(n21137), .B2(
        gray_img[31]), .O(n21809) );
  AOI22S U27370 ( .A1(n22920), .A2(gray_img[663]), .B1(gray_img[919]), .B2(
        n22894), .O(n21808) );
  AOI22S U27371 ( .A1(n22895), .A2(gray_img[407]), .B1(gray_img[1687]), .B2(
        n22896), .O(n21807) );
  ND3S U27372 ( .I1(n21809), .I2(n21808), .I3(n21807), .O(n21821) );
  AOI22S U27373 ( .A1(n15921), .A2(gray_img[1175]), .B1(gray_img[1559]), .B2(
        n15919), .O(n21819) );
  ND2S U27374 ( .I1(n22819), .I2(gray_img[927]), .O(n21816) );
  ND2S U27375 ( .I1(n22900), .I2(gray_img[15]), .O(n21815) );
  ND2S U27376 ( .I1(n22812), .I2(gray_img[1927]), .O(n21814) );
  AOI22S U27377 ( .A1(gray_img[159]), .A2(n21089), .B1(gray_img[535]), .B2(
        n15915), .O(n21812) );
  AOI22S U27378 ( .A1(gray_img[23]), .A2(n22901), .B1(gray_img[1943]), .B2(
        n22679), .O(n21811) );
  ND2S U27379 ( .I1(gray_img[1047]), .I2(n22929), .O(n21810) );
  ND3S U27380 ( .I1(n21812), .I2(n21811), .I3(n21810), .O(n21813) );
  AN4B1S U27381 ( .I1(n21816), .I2(n21815), .I3(n21814), .B1(n21813), .O(
        n21818) );
  AOI22S U27382 ( .A1(n22566), .A2(gray_img[903]), .B1(gray_img[391]), .B2(
        n22686), .O(n21817) );
  ND3S U27383 ( .I1(n21819), .I2(n21818), .I3(n21817), .O(n21820) );
  AO112S U27384 ( .C1(gray_img[7]), .C2(n22893), .A1(n21821), .B1(n21820), .O(
        n21822) );
  NR3 U27385 ( .I1(n21824), .I2(n21823), .I3(n21822), .O(n21825) );
  ND3S U27386 ( .I1(n21827), .I2(n21826), .I3(n21825), .O(n21883) );
  AOI22S U27387 ( .A1(n22727), .A2(gray_img[1903]), .B1(n22895), .B2(
        gray_img[503]), .O(n21832) );
  AOI22S U27388 ( .A1(n22810), .A2(gray_img[743]), .B1(gray_img[1007]), .B2(
        n22802), .O(n21831) );
  AOI22S U27389 ( .A1(n22657), .A2(gray_img[751]), .B1(gray_img[1791]), .B2(
        n22505), .O(n21830) );
  MOAI1S U27390 ( .A1(n21828), .A2(n27568), .B1(n22867), .B2(gray_img[895]), 
        .O(n21829) );
  AN4B1S U27391 ( .I1(n21832), .I2(n21831), .I3(n21830), .B1(n21829), .O(
        n21881) );
  AOI22S U27392 ( .A1(n22921), .A2(gray_img[1775]), .B1(gray_img[1263]), .B2(
        n22936), .O(n21836) );
  AOI22S U27393 ( .A1(n22837), .A2(gray_img[367]), .B1(gray_img[1127]), .B2(
        n22703), .O(n21835) );
  AOI22S U27394 ( .A1(n22630), .A2(gray_img[615]), .B1(gray_img[511]), .B2(
        n22881), .O(n21834) );
  MOAI1S U27395 ( .A1(n25792), .A2(n22218), .B1(n22664), .B2(gray_img[1527]), 
        .O(n21833) );
  AN4B1S U27396 ( .I1(n21836), .I2(n21835), .I3(n21834), .B1(n21833), .O(
        n21880) );
  AOI22S U27397 ( .A1(n22735), .A2(gray_img[383]), .B1(gray_img[1511]), .B2(
        n21106), .O(n21840) );
  ND2S U27398 ( .I1(n22863), .I2(gray_img[1911]), .O(n21839) );
  AOI22S U27399 ( .A1(n22887), .A2(gray_img[623]), .B1(gray_img[767]), .B2(
        n22883), .O(n21838) );
  INV1S U27400 ( .I(gray_img[1639]), .O(n25804) );
  MOAI1S U27401 ( .A1(n22670), .A2(n25804), .B1(n22872), .B2(gray_img[1255]), 
        .O(n21837) );
  AN4B1S U27402 ( .I1(n21840), .I2(n21839), .I3(n21838), .B1(n21837), .O(
        n21859) );
  INV1S U27403 ( .I(gray_img[999]), .O(n26255) );
  MOAI1S U27404 ( .A1(n21841), .A2(n26255), .B1(n22686), .B2(gray_img[487]), 
        .O(n21852) );
  INV1S U27405 ( .I(gray_img[1399]), .O(n27917) );
  NR2 U27406 ( .I1(n27917), .I2(n22797), .O(n21851) );
  ND2S U27407 ( .I1(n22827), .I2(gray_img[1655]), .O(n21849) );
  ND2S U27408 ( .I1(n22900), .I2(gray_img[111]), .O(n21846) );
  AOI22S U27409 ( .A1(gray_img[119]), .A2(n22901), .B1(gray_img[1663]), .B2(
        n22918), .O(n21845) );
  ND2S U27410 ( .I1(n22812), .I2(gray_img[2023]), .O(n21844) );
  INV1S U27411 ( .I(gray_img[1143]), .O(n23311) );
  MOAI1S U27412 ( .A1(n23311), .A2(n21842), .B1(gray_img[2039]), .B2(n22679), 
        .O(n21843) );
  AN4B1S U27413 ( .I1(n21846), .I2(n21845), .I3(n21844), .B1(n21843), .O(
        n21848) );
  ND2S U27414 ( .I1(n22819), .I2(gray_img[1023]), .O(n21847) );
  ND3S U27415 ( .I1(n21849), .I2(n21848), .I3(n21847), .O(n21850) );
  NR3 U27416 ( .I1(n21852), .I2(n21851), .I3(n21850), .O(n21858) );
  ND2S U27417 ( .I1(n22893), .I2(gray_img[103]), .O(n21857) );
  ND2S U27418 ( .I1(n15918), .I2(gray_img[247]), .O(n21855) );
  AOI22S U27419 ( .A1(n22770), .A2(gray_img[1767]), .B1(gray_img[359]), .B2(
        n22625), .O(n21854) );
  AOI22S U27420 ( .A1(n22513), .A2(gray_img[871]), .B1(gray_img[231]), .B2(
        n22610), .O(n21853) );
  ND3S U27421 ( .I1(n21855), .I2(n21854), .I3(n21853), .O(n21856) );
  AN4B1S U27422 ( .I1(n21859), .I2(n21858), .I3(n21857), .B1(n21856), .O(
        n21866) );
  AOI22S U27423 ( .A1(n21096), .A2(gray_img[1535]), .B1(gray_img[1279]), .B2(
        n21090), .O(n21865) );
  ND2S U27424 ( .I1(n22755), .I2(gray_img[2047]), .O(n21864) );
  AOI22S U27425 ( .A1(n21120), .A2(gray_img[1407]), .B1(n21137), .B2(
        gray_img[127]), .O(n21862) );
  AOI22S U27426 ( .A1(n22695), .A2(gray_img[759]), .B1(gray_img[1015]), .B2(
        n22894), .O(n21861) );
  AOI22S U27427 ( .A1(n22896), .A2(gray_img[1783]), .B1(gray_img[1271]), .B2(
        n15921), .O(n21860) );
  ND3S U27428 ( .I1(n21862), .I2(n21861), .I3(n21860), .O(n21863) );
  AN4B1S U27429 ( .I1(n21866), .I2(n21865), .I3(n21864), .B1(n21863), .O(
        n21878) );
  AOI22S U27430 ( .A1(n15905), .A2(gray_img[375]), .B1(gray_img[887]), .B2(
        n22930), .O(n21877) );
  ND2S U27431 ( .I1(n21152), .I2(gray_img[639]), .O(n21870) );
  AOI22S U27432 ( .A1(n22794), .A2(gray_img[1895]), .B1(gray_img[1135]), .B2(
        n21155), .O(n21869) );
  AOI22S U27433 ( .A1(n22787), .A2(gray_img[1919]), .B1(gray_img[1383]), .B2(
        n22934), .O(n21868) );
  MOAI1S U27434 ( .A1(n22875), .A2(n27984), .B1(n22861), .B2(gray_img[1391]), 
        .O(n21867) );
  AN4B1S U27435 ( .I1(n21870), .I2(n21869), .I3(n21868), .B1(n21867), .O(
        n21871) );
  OA12S U27436 ( .B1(n25860), .B2(n22853), .A1(n21871), .O(n21876) );
  ND2S U27437 ( .I1(n15915), .I2(gray_img[631]), .O(n21874) );
  AOI22S U27438 ( .A1(n22933), .A2(gray_img[239]), .B1(gray_img[879]), .B2(
        n22724), .O(n21873) );
  AOI22S U27439 ( .A1(n22762), .A2(gray_img[495]), .B1(gray_img[1151]), .B2(
        n22935), .O(n21872) );
  ND3S U27440 ( .I1(n21874), .I2(n21873), .I3(n21872), .O(n21875) );
  AN4B1S U27441 ( .I1(n21878), .I2(n21877), .I3(n21876), .B1(n21875), .O(
        n21879) );
  AOI22S U27442 ( .A1(n22784), .A2(n21883), .B1(n22959), .B2(n21882), .O(
        n21988) );
  INV1S U27443 ( .I(gray_img[719]), .O(n27158) );
  MOAI1S U27444 ( .A1(n21884), .A2(n27158), .B1(n22785), .B2(gray_img[351]), 
        .O(n21890) );
  MOAI1S U27445 ( .A1(n22218), .A2(n25666), .B1(n22836), .B2(gray_img[207]), 
        .O(n21889) );
  ND2S U27446 ( .I1(n21096), .I2(gray_img[1503]), .O(n21887) );
  AOI22S U27447 ( .A1(gray_img[223]), .A2(n21089), .B1(n22819), .B2(
        gray_img[991]), .O(n21886) );
  ND2S U27448 ( .I1(n15921), .I2(gray_img[1239]), .O(n21885) );
  ND3S U27449 ( .I1(n21887), .I2(n21886), .I3(n21885), .O(n21888) );
  NR3 U27450 ( .I1(n21890), .I2(n21889), .I3(n21888), .O(n21932) );
  AOI22S U27451 ( .A1(n22921), .A2(gray_img[1743]), .B1(n22796), .B2(
        gray_img[1751]), .O(n21894) );
  AOI22S U27452 ( .A1(gray_img[607]), .A2(n21152), .B1(n22630), .B2(
        gray_img[583]), .O(n21893) );
  AOI22S U27453 ( .A1(n22770), .A2(gray_img[1735]), .B1(gray_img[327]), .B2(
        n22625), .O(n21892) );
  MOAI1S U27454 ( .A1(n22346), .A2(n22982), .B1(n22686), .B2(gray_img[455]), 
        .O(n21891) );
  AN4B1S U27455 ( .I1(n21894), .I2(n21893), .I3(n21892), .B1(n21891), .O(
        n21931) );
  AOI22S U27456 ( .A1(n22863), .A2(gray_img[1879]), .B1(gray_img[1367]), .B2(
        n22889), .O(n21900) );
  AOI22S U27457 ( .A1(n22909), .A2(gray_img[711]), .B1(gray_img[591]), .B2(
        n22795), .O(n21899) );
  ND2S U27458 ( .I1(n22911), .I2(gray_img[967]), .O(n21898) );
  INV1S U27459 ( .I(gray_img[79]), .O(n23601) );
  AOI22S U27460 ( .A1(gray_img[2007]), .A2(n22679), .B1(gray_img[87]), .B2(
        n22901), .O(n21896) );
  ND2S U27461 ( .I1(n22812), .I2(gray_img[1991]), .O(n21895) );
  OAI112HS U27462 ( .C1(n22811), .C2(n23601), .A1(n21896), .B1(n21895), .O(
        n21897) );
  AN4B1S U27463 ( .I1(n21900), .I2(n21899), .I3(n21898), .B1(n21897), .O(
        n21908) );
  AOI22S U27464 ( .A1(n22881), .A2(gray_img[479]), .B1(gray_img[1607]), .B2(
        n21097), .O(n21904) );
  AOI22S U27465 ( .A1(n22513), .A2(gray_img[839]), .B1(gray_img[199]), .B2(
        n22610), .O(n21903) );
  AOI22S U27466 ( .A1(n22505), .A2(gray_img[1759]), .B1(gray_img[735]), .B2(
        n22883), .O(n21902) );
  INV1S U27467 ( .I(gray_img[1479]), .O(n23511) );
  MOAI1S U27468 ( .A1(n22718), .A2(n23511), .B1(n22872), .B2(gray_img[1223]), 
        .O(n21901) );
  AN4B1S U27469 ( .I1(n21904), .I2(n21903), .I3(n21902), .B1(n21901), .O(
        n21907) );
  AOI22S U27470 ( .A1(n15918), .A2(gray_img[215]), .B1(gray_img[343]), .B2(
        n15905), .O(n21906) );
  INV1S U27471 ( .I(gray_img[855]), .O(n23066) );
  MOAI1S U27472 ( .A1(n22841), .A2(n23066), .B1(n15915), .B2(gray_img[599]), 
        .O(n21905) );
  AN4B1S U27473 ( .I1(n21908), .I2(n21907), .I3(n21906), .B1(n21905), .O(
        n21929) );
  ND2S U27474 ( .I1(n22929), .I2(gray_img[1111]), .O(n21912) );
  AOI22S U27475 ( .A1(n22837), .A2(gray_img[335]), .B1(gray_img[847]), .B2(
        n22932), .O(n21911) );
  AOI22S U27476 ( .A1(n22762), .A2(gray_img[463]), .B1(gray_img[1119]), .B2(
        n22935), .O(n21910) );
  NR2 U27477 ( .I1(n25001), .I2(n22853), .O(n21909) );
  AN4B1S U27478 ( .I1(n21912), .I2(n21911), .I3(n21910), .B1(n21909), .O(
        n21928) );
  AOI22S U27479 ( .A1(n22695), .A2(gray_img[727]), .B1(gray_img[983]), .B2(
        n22894), .O(n21918) );
  AOI22S U27480 ( .A1(n22664), .A2(gray_img[1495]), .B1(gray_img[1623]), .B2(
        n15919), .O(n21917) );
  ND2S U27481 ( .I1(n22893), .I2(gray_img[71]), .O(n21916) );
  ND2S U27482 ( .I1(n22919), .I2(gray_img[2015]), .O(n21914) );
  AOI22S U27483 ( .A1(n22937), .A2(gray_img[1871]), .B1(n22895), .B2(
        gray_img[471]), .O(n21913) );
  OAI112HS U27484 ( .C1(n22924), .C2(n25222), .A1(n21914), .B1(n21913), .O(
        n21915) );
  AN4B1S U27485 ( .I1(n21918), .I2(n21917), .I3(n21916), .B1(n21915), .O(
        n21927) );
  AOI22S U27486 ( .A1(n21155), .A2(gray_img[1103]), .B1(gray_img[1231]), .B2(
        n22936), .O(n21922) );
  AOI22S U27487 ( .A1(n22934), .A2(gray_img[1351]), .B1(gray_img[1095]), .B2(
        n22703), .O(n21921) );
  AOI22S U27488 ( .A1(n22787), .A2(gray_img[1887]), .B1(gray_img[1863]), .B2(
        n22938), .O(n21920) );
  INV1S U27489 ( .I(gray_img[1487]), .O(n25199) );
  MOAI1S U27490 ( .A1(n22875), .A2(n25199), .B1(n22861), .B2(gray_img[1359]), 
        .O(n21919) );
  AN4B1S U27491 ( .I1(n21922), .I2(n21921), .I3(n21920), .B1(n21919), .O(
        n21925) );
  AOI22S U27492 ( .A1(n22867), .A2(gray_img[863]), .B1(gray_img[1631]), .B2(
        n22694), .O(n21924) );
  AOI22S U27493 ( .A1(n21090), .A2(gray_img[1247]), .B1(gray_img[1375]), .B2(
        n21120), .O(n21923) );
  AN4B1S U27494 ( .I1(n21929), .I2(n21928), .I3(n21927), .B1(n21926), .O(
        n21930) );
  ND3S U27495 ( .I1(n21932), .I2(n21931), .I3(n21930), .O(n21986) );
  MOAI1S U27496 ( .A1(n21933), .A2(n28169), .B1(n22895), .B2(gray_img[439]), 
        .O(n21940) );
  NR2 U27497 ( .I1(n21934), .I2(n22493), .O(n21939) );
  AOI22S U27498 ( .A1(n22896), .A2(gray_img[1719]), .B1(gray_img[1591]), .B2(
        n15919), .O(n21937) );
  AOI22S U27499 ( .A1(n22610), .A2(gray_img[167]), .B1(gray_img[815]), .B2(
        n22932), .O(n21936) );
  ND2S U27500 ( .I1(n22867), .I2(gray_img[831]), .O(n21935) );
  ND3S U27501 ( .I1(n21937), .I2(n21936), .I3(n21935), .O(n21938) );
  NR3 U27502 ( .I1(n21940), .I2(n21939), .I3(n21938), .O(n21984) );
  AOI22S U27503 ( .A1(n22938), .A2(gray_img[1831]), .B1(n22664), .B2(
        gray_img[1463]), .O(n21944) );
  AOI22S U27504 ( .A1(n22836), .A2(gray_img[175]), .B1(gray_img[431]), .B2(
        n22762), .O(n21943) );
  AOI22S U27505 ( .A1(n22795), .A2(gray_img[559]), .B1(gray_img[295]), .B2(
        n22625), .O(n21942) );
  INV1S U27506 ( .I(gray_img[1207]), .O(n28878) );
  MOAI1S U27507 ( .A1(n28878), .A2(n22058), .B1(n22889), .B2(gray_img[1335]), 
        .O(n21941) );
  AN4B1S U27508 ( .I1(n21944), .I2(n21943), .I3(n21942), .B1(n21941), .O(
        n21983) );
  AOI22S U27509 ( .A1(n22910), .A2(gray_img[943]), .B1(gray_img[687]), .B2(
        n22888), .O(n21948) );
  ND2S U27510 ( .I1(n22863), .I2(gray_img[1847]), .O(n21947) );
  AOI22S U27511 ( .A1(n22911), .A2(gray_img[935]), .B1(gray_img[679]), .B2(
        n22909), .O(n21946) );
  INV1S U27512 ( .I(gray_img[1727]), .O(n29209) );
  MOAI1S U27513 ( .A1(n22882), .A2(n29209), .B1(n22883), .B2(gray_img[703]), 
        .O(n21945) );
  AN4B1S U27514 ( .I1(n21948), .I2(n21947), .I3(n21946), .B1(n21945), .O(
        n21956) );
  AOI22S U27515 ( .A1(n21155), .A2(gray_img[1071]), .B1(n22828), .B2(
        gray_img[951]), .O(n21955) );
  AOI22S U27516 ( .A1(n22630), .A2(gray_img[551]), .B1(gray_img[423]), .B2(
        n22686), .O(n21954) );
  INV1S U27517 ( .I(gray_img[47]), .O(n26968) );
  ND2S U27518 ( .I1(n22819), .I2(gray_img[959]), .O(n21952) );
  AOI22S U27519 ( .A1(gray_img[55]), .A2(n22901), .B1(gray_img[1215]), .B2(
        n21090), .O(n21950) );
  ND2S U27520 ( .I1(gray_img[1975]), .I2(n22679), .O(n21949) );
  OAI112HS U27521 ( .C1(n22811), .C2(n26968), .A1(n21952), .B1(n21951), .O(
        n21953) );
  AN4B1S U27522 ( .I1(n21956), .I2(n21955), .I3(n21954), .B1(n21953), .O(
        n21981) );
  AOI22S U27523 ( .A1(n21120), .A2(gray_img[1343]), .B1(n21137), .B2(
        gray_img[63]), .O(n21960) );
  AOI22S U27524 ( .A1(n21089), .A2(gray_img[191]), .B1(gray_img[1599]), .B2(
        n22694), .O(n21959) );
  ND2S U27525 ( .I1(n22893), .I2(gray_img[39]), .O(n21958) );
  INV1S U27526 ( .I(gray_img[1983]), .O(n23138) );
  NR2 U27527 ( .I1(n23138), .I2(n22251), .O(n21957) );
  AN4B1S U27528 ( .I1(n21960), .I2(n21959), .I3(n21958), .B1(n21957), .O(
        n21980) );
  AOI22S U27529 ( .A1(n22785), .A2(gray_img[319]), .B1(gray_img[447]), .B2(
        n22881), .O(n21964) );
  AOI22S U27530 ( .A1(n21106), .A2(gray_img[1447]), .B1(gray_img[1575]), .B2(
        n21097), .O(n21963) );
  ND2S U27531 ( .I1(n15918), .I2(gray_img[183]), .O(n21962) );
  INV1S U27532 ( .I(gray_img[311]), .O(n26513) );
  MOAI1S U27533 ( .A1(n22383), .A2(n26513), .B1(n22930), .B2(gray_img[823]), 
        .O(n21961) );
  AN4B1S U27534 ( .I1(n21964), .I2(n21963), .I3(n21962), .B1(n21961), .O(
        n21979) );
  ND2S U27535 ( .I1(n22929), .I2(gray_img[1079]), .O(n21971) );
  AOI22S U27536 ( .A1(n22935), .A2(gray_img[1087]), .B1(gray_img[1855]), .B2(
        n22787), .O(n21970) );
  AOI22S U27537 ( .A1(n22934), .A2(gray_img[1319]), .B1(gray_img[1063]), .B2(
        n22703), .O(n21969) );
  ND2S U27538 ( .I1(n15915), .I2(gray_img[567]), .O(n21967) );
  AOI22S U27539 ( .A1(n22770), .A2(gray_img[1703]), .B1(gray_img[1191]), .B2(
        n22838), .O(n21966) );
  AOI22S U27540 ( .A1(n22513), .A2(gray_img[807]), .B1(gray_img[303]), .B2(
        n22837), .O(n21965) );
  ND3S U27541 ( .I1(n21967), .I2(n21966), .I3(n21965), .O(n21968) );
  AN4B1S U27542 ( .I1(n21971), .I2(n21970), .I3(n21969), .B1(n21968), .O(
        n21977) );
  AOI22S U27543 ( .A1(n22656), .A2(gray_img[1583]), .B1(gray_img[1455]), .B2(
        n22369), .O(n21975) );
  AOI22S U27544 ( .A1(n22846), .A2(gray_img[1327]), .B1(gray_img[1711]), .B2(
        n22921), .O(n21974) );
  AOI22S U27545 ( .A1(n22937), .A2(gray_img[1839]), .B1(gray_img[1199]), .B2(
        n22936), .O(n21973) );
  INV1S U27546 ( .I(gray_img[575]), .O(n28154) );
  NR2 U27547 ( .I1(n28154), .I2(n22750), .O(n21972) );
  AN4B1S U27548 ( .I1(n21975), .I2(n21974), .I3(n21973), .B1(n21972), .O(
        n21976) );
  OAI112HS U27549 ( .C1(n26681), .C2(n22853), .A1(n21977), .B1(n21976), .O(
        n21978) );
  AN4B1S U27550 ( .I1(n21981), .I2(n21980), .I3(n21979), .B1(n21978), .O(
        n21982) );
  AOI22S U27551 ( .A1(n22782), .A2(n21986), .B1(n22957), .B2(n21985), .O(
        n21987) );
  ND2S U27552 ( .I1(n21089), .I2(gray_img[216]), .O(n21994) );
  AOI22S U27553 ( .A1(n22610), .A2(gray_img[192]), .B1(gray_img[200]), .B2(
        n22836), .O(n21993) );
  AOI22S U27554 ( .A1(n22630), .A2(gray_img[576]), .B1(gray_img[472]), .B2(
        n22881), .O(n21992) );
  ND2S U27555 ( .I1(n22828), .I2(gray_img[976]), .O(n21990) );
  AOI22S U27556 ( .A1(gray_img[1624]), .A2(n22918), .B1(n22566), .B2(
        gray_img[960]), .O(n21989) );
  ND2S U27557 ( .I1(n21990), .I2(n21989), .O(n21991) );
  AN4B1S U27558 ( .I1(n21994), .I2(n21993), .I3(n21992), .B1(n21991), .O(
        n22045) );
  ND2S U27559 ( .I1(n22930), .I2(gray_img[848]), .O(n22001) );
  AOI22S U27560 ( .A1(n22770), .A2(gray_img[1728]), .B1(gray_img[456]), .B2(
        n22762), .O(n22000) );
  ND2S U27561 ( .I1(n21152), .I2(gray_img[600]), .O(n21999) );
  ND2S U27562 ( .I1(n21096), .I2(gray_img[1496]), .O(n21997) );
  AOI22S U27563 ( .A1(n22887), .A2(gray_img[584]), .B1(gray_img[344]), .B2(
        n22785), .O(n21996) );
  ND2S U27564 ( .I1(n21155), .I2(gray_img[1096]), .O(n21995) );
  ND3S U27565 ( .I1(n21997), .I2(n21996), .I3(n21995), .O(n21998) );
  AN4B1S U27566 ( .I1(n22001), .I2(n22000), .I3(n21999), .B1(n21998), .O(
        n22044) );
  ND2S U27567 ( .I1(n22893), .I2(gray_img[64]), .O(n22014) );
  AOI22S U27568 ( .A1(n22802), .A2(gray_img[968]), .B1(gray_img[712]), .B2(
        n22888), .O(n22013) );
  ND2S U27569 ( .I1(n22863), .I2(gray_img[1872]), .O(n22012) );
  AOI22S U27570 ( .A1(n22810), .A2(gray_img[704]), .B1(gray_img[448]), .B2(
        n22686), .O(n22010) );
  AOI22S U27571 ( .A1(gray_img[856]), .A2(n22813), .B1(gray_img[1240]), .B2(
        n21090), .O(n22004) );
  AOI22S U27572 ( .A1(gray_img[1104]), .A2(n22929), .B1(gray_img[2000]), .B2(
        n22679), .O(n22003) );
  ND2S U27573 ( .I1(gray_img[80]), .I2(n22901), .O(n22002) );
  ND3S U27574 ( .I1(n22004), .I2(n22003), .I3(n22002), .O(n22007) );
  NR2 U27575 ( .I1(intadd_130_A_0_), .I2(n22811), .O(n22006) );
  NR2 U27576 ( .I1(intadd_25_A_0_), .I2(n22904), .O(n22005) );
  NR3 U27577 ( .I1(n22007), .I2(n22006), .I3(n22005), .O(n22009) );
  ND2S U27578 ( .I1(n22819), .I2(gray_img[984]), .O(n22008) );
  AN4B1S U27579 ( .I1(n22014), .I2(n22013), .I3(n22012), .B1(n22011), .O(
        n22019) );
  AOI22S U27580 ( .A1(n22796), .A2(gray_img[1744]), .B1(gray_img[1616]), .B2(
        n15919), .O(n22018) );
  AOI22S U27581 ( .A1(n22664), .A2(gray_img[1488]), .B1(gray_img[1232]), .B2(
        n15921), .O(n22017) );
  AOI22S U27582 ( .A1(n22895), .A2(gray_img[464]), .B1(gray_img[720]), .B2(
        n22920), .O(n22015) );
  OAI12HS U27583 ( .B1(n22924), .B2(intadd_188_A_0_), .A1(n22015), .O(n22016)
         );
  AN4B1S U27584 ( .I1(n22019), .I2(n22018), .I3(n22017), .B1(n22016), .O(
        n22042) );
  ND2S U27585 ( .I1(n22931), .I2(gray_img[1992]), .O(n22030) );
  AOI22S U27586 ( .A1(n22786), .A2(gray_img[1752]), .B1(gray_img[728]), .B2(
        n22883), .O(n22023) );
  AOI22S U27587 ( .A1(n22872), .A2(gray_img[1216]), .B1(gray_img[320]), .B2(
        n22625), .O(n22022) );
  ND2S U27588 ( .I1(n22889), .I2(gray_img[1360]), .O(n22021) );
  MOAI1S U27589 ( .A1(n22718), .A2(intadd_186_A_0_), .B1(n21097), .B2(
        gray_img[1600]), .O(n22020) );
  AN4B1S U27590 ( .I1(n22023), .I2(n22022), .I3(n22021), .B1(n22020), .O(
        n22029) );
  AOI22S U27591 ( .A1(n15918), .A2(gray_img[208]), .B1(gray_img[336]), .B2(
        n15905), .O(n22028) );
  ND2S U27592 ( .I1(n15915), .I2(gray_img[592]), .O(n22026) );
  AOI22S U27593 ( .A1(n22513), .A2(gray_img[832]), .B1(gray_img[840]), .B2(
        n22932), .O(n22025) );
  AOI22S U27594 ( .A1(n22837), .A2(gray_img[328]), .B1(gray_img[1112]), .B2(
        n22935), .O(n22024) );
  ND3S U27595 ( .I1(n22026), .I2(n22025), .I3(n22024), .O(n22027) );
  AN4B1S U27596 ( .I1(n22030), .I2(n22029), .I3(n22028), .B1(n22027), .O(
        n22041) );
  AOI22S U27597 ( .A1(n22921), .A2(gray_img[1736]), .B1(gray_img[1224]), .B2(
        n22936), .O(n22035) );
  AOI22S U27598 ( .A1(n22934), .A2(gray_img[1344]), .B1(gray_img[1088]), .B2(
        n22703), .O(n22034) );
  AOI22S U27599 ( .A1(n22787), .A2(gray_img[1880]), .B1(gray_img[1856]), .B2(
        n22794), .O(n22033) );
  MOAI1S U27600 ( .A1(n22031), .A2(n30458), .B1(n22727), .B2(gray_img[1864]), 
        .O(n22032) );
  AN4B1S U27601 ( .I1(n22035), .I2(n22034), .I3(n22033), .B1(n22032), .O(
        n22040) );
  ND2S U27602 ( .I1(n22919), .I2(gray_img[2008]), .O(n22038) );
  AOI22S U27603 ( .A1(n22874), .A2(gray_img[1608]), .B1(gray_img[1480]), .B2(
        n22369), .O(n22037) );
  ND2S U27604 ( .I1(n21120), .I2(gray_img[1368]), .O(n22036) );
  ND3S U27605 ( .I1(n22038), .I2(n22037), .I3(n22036), .O(n22039) );
  AN4B1S U27606 ( .I1(n22042), .I2(n22041), .I3(n22040), .B1(n22039), .O(
        n22043) );
  AOI22S U27607 ( .A1(n22921), .A2(gray_img[1704]), .B1(n22664), .B2(
        gray_img[1456]), .O(n22050) );
  AOI22S U27608 ( .A1(n22883), .A2(gray_img[696]), .B1(gray_img[1184]), .B2(
        n22872), .O(n22049) );
  AOI22S U27609 ( .A1(n21106), .A2(gray_img[1440]), .B1(n22703), .B2(
        gray_img[1056]), .O(n22048) );
  MOAI1S U27610 ( .A1(n22156), .A2(n22046), .B1(n22911), .B2(gray_img[928]), 
        .O(n22047) );
  AN4B1S U27611 ( .I1(n22050), .I2(n22049), .I3(n22048), .B1(n22047), .O(
        n22099) );
  AOI22S U27612 ( .A1(n22938), .A2(gray_img[1824]), .B1(gray_img[1320]), .B2(
        n22861), .O(n22056) );
  AOI22S U27613 ( .A1(n22686), .A2(gray_img[416]), .B1(gray_img[680]), .B2(
        n22657), .O(n22055) );
  ND2S U27614 ( .I1(n21155), .I2(gray_img[1064]), .O(n22054) );
  AOI22S U27615 ( .A1(n22724), .A2(gray_img[808]), .B1(gray_img[1312]), .B2(
        n22934), .O(n22052) );
  ND2S U27616 ( .I1(n22863), .I2(gray_img[1840]), .O(n22051) );
  ND2S U27617 ( .I1(n22052), .I2(n22051), .O(n22053) );
  AN4B1S U27618 ( .I1(n22056), .I2(n22055), .I3(n22054), .B1(n22053), .O(
        n22098) );
  AOI22S U27619 ( .A1(n22619), .A2(gray_img[432]), .B1(gray_img[944]), .B2(
        n22894), .O(n22062) );
  AOI22S U27620 ( .A1(n22920), .A2(gray_img[688]), .B1(gray_img[1584]), .B2(
        n15919), .O(n22061) );
  ND2S U27621 ( .I1(n21137), .I2(gray_img[56]), .O(n22060) );
  INV1S U27622 ( .I(gray_img[1200]), .O(n22057) );
  MOAI1S U27623 ( .A1(n22058), .A2(n22057), .B1(n22796), .B2(gray_img[1712]), 
        .O(n22059) );
  AN4B1S U27624 ( .I1(n22062), .I2(n22061), .I3(n22060), .B1(n22059), .O(
        n22065) );
  AOI22S U27625 ( .A1(n21090), .A2(gray_img[1208]), .B1(gray_img[1336]), .B2(
        n21120), .O(n22064) );
  ND2S U27626 ( .I1(n22755), .I2(gray_img[1976]), .O(n22063) );
  AOI22S U27627 ( .A1(n22735), .A2(gray_img[312]), .B1(gray_img[440]), .B2(
        n22736), .O(n22069) );
  AOI22S U27628 ( .A1(n22770), .A2(gray_img[1696]), .B1(gray_img[1568]), .B2(
        n21097), .O(n22068) );
  ND2S U27629 ( .I1(n15918), .I2(gray_img[176]), .O(n22067) );
  MOAI1S U27630 ( .A1(n22841), .A2(n26097), .B1(n15915), .B2(gray_img[560]), 
        .O(n22066) );
  AN4B1S U27631 ( .I1(n22069), .I2(n22068), .I3(n22067), .B1(n22066), .O(
        n22081) );
  AOI22S U27632 ( .A1(n22887), .A2(gray_img[552]), .B1(gray_img[1720]), .B2(
        n22505), .O(n22078) );
  ND2S U27633 ( .I1(n22889), .I2(gray_img[1328]), .O(n22077) );
  AOI22S U27634 ( .A1(n22630), .A2(gray_img[544]), .B1(gray_img[936]), .B2(
        n22910), .O(n22076) );
  ND2S U27635 ( .I1(n22819), .I2(gray_img[952]), .O(n22074) );
  INV1S U27636 ( .I(gray_img[40]), .O(n26956) );
  AOI22S U27637 ( .A1(gray_img[48]), .A2(n22901), .B1(gray_img[304]), .B2(
        n15905), .O(n22071) );
  AOI22S U27638 ( .A1(gray_img[1968]), .A2(n22679), .B1(gray_img[1464]), .B2(
        n21096), .O(n22070) );
  OA112S U27639 ( .C1(n22811), .C2(n26956), .A1(n22071), .B1(n22070), .O(
        n22073) );
  ND2S U27640 ( .I1(n22812), .I2(gray_img[1952]), .O(n22072) );
  ND3S U27641 ( .I1(n22074), .I2(n22073), .I3(n22072), .O(n22075) );
  AN4B1S U27642 ( .I1(n22078), .I2(n22077), .I3(n22076), .B1(n22075), .O(
        n22080) );
  ND2S U27643 ( .I1(n22893), .I2(gray_img[32]), .O(n22079) );
  ND3S U27644 ( .I1(n22081), .I2(n22080), .I3(n22079), .O(n22095) );
  AOI22S U27645 ( .A1(n22874), .A2(gray_img[1576]), .B1(gray_img[1448]), .B2(
        n22369), .O(n22085) );
  AOI22S U27646 ( .A1(n22727), .A2(gray_img[1832]), .B1(gray_img[1192]), .B2(
        n22936), .O(n22084) );
  AOI22S U27647 ( .A1(n22935), .A2(gray_img[1080]), .B1(gray_img[1848]), .B2(
        n22864), .O(n22083) );
  MOAI1S U27648 ( .A1(n22865), .A2(intadd_16_B_0_), .B1(n22933), .B2(
        gray_img[168]), .O(n22082) );
  AN4B1S U27649 ( .I1(n22085), .I2(n22084), .I3(n22083), .B1(n22082), .O(
        n22088) );
  AOI22S U27650 ( .A1(n21152), .A2(gray_img[568]), .B1(gray_img[824]), .B2(
        n22813), .O(n22087) );
  AOI22S U27651 ( .A1(n21089), .A2(gray_img[184]), .B1(gray_img[1592]), .B2(
        n22694), .O(n22086) );
  ND3S U27652 ( .I1(n22088), .I2(n22087), .I3(n22086), .O(n22093) );
  ND2S U27653 ( .I1(n22929), .I2(gray_img[1072]), .O(n22091) );
  AOI22S U27654 ( .A1(n22513), .A2(gray_img[800]), .B1(gray_img[160]), .B2(
        n22610), .O(n22090) );
  AOI22S U27655 ( .A1(n22625), .A2(gray_img[288]), .B1(gray_img[424]), .B2(
        n22762), .O(n22089) );
  ND3S U27656 ( .I1(n22091), .I2(n22090), .I3(n22089), .O(n22092) );
  AO112S U27657 ( .C1(gray_img[1960]), .C2(n22931), .A1(n22093), .B1(n22092), 
        .O(n22094) );
  NR3 U27658 ( .I1(n22096), .I2(n22095), .I3(n22094), .O(n22097) );
  ND3S U27659 ( .I1(n22099), .I2(n22098), .I3(n22097), .O(n22100) );
  AOI22S U27660 ( .A1(n22782), .A2(n22101), .B1(n22957), .B2(n22100), .O(
        n22217) );
  AOI22S U27661 ( .A1(n15921), .A2(gray_img[1168]), .B1(gray_img[1552]), .B2(
        n15919), .O(n22107) );
  AOI22S U27662 ( .A1(n22881), .A2(gray_img[408]), .B1(gray_img[1536]), .B2(
        n21097), .O(n22106) );
  AOI22S U27663 ( .A1(n22703), .A2(gray_img[1024]), .B1(gray_img[1160]), .B2(
        n22936), .O(n22105) );
  MOAI1S U27664 ( .A1(n22103), .A2(n22102), .B1(n22657), .B2(gray_img[648]), 
        .O(n22104) );
  AN4B1S U27665 ( .I1(n22107), .I2(n22106), .I3(n22105), .B1(n22104), .O(
        n22155) );
  AOI22S U27666 ( .A1(n22762), .A2(gray_img[392]), .B1(n22921), .B2(
        gray_img[1672]), .O(n22112) );
  AOI22S U27667 ( .A1(n22802), .A2(gray_img[904]), .B1(gray_img[520]), .B2(
        n22795), .O(n22111) );
  AOI22S U27668 ( .A1(n22873), .A2(gray_img[920]), .B1(gray_img[384]), .B2(
        n22686), .O(n22110) );
  INV1S U27669 ( .I(gray_img[1152]), .O(n22108) );
  MOAI1S U27670 ( .A1(n22392), .A2(n22108), .B1(n22505), .B2(gray_img[1688]), 
        .O(n22109) );
  AN4B1S U27671 ( .I1(n22112), .I2(n22111), .I3(n22110), .B1(n22109), .O(
        n22154) );
  AOI22S U27672 ( .A1(n15918), .A2(gray_img[144]), .B1(gray_img[272]), .B2(
        n15905), .O(n22116) );
  AOI22S U27673 ( .A1(n22883), .A2(gray_img[664]), .B1(gray_img[280]), .B2(
        n22735), .O(n22115) );
  AOI22S U27674 ( .A1(n21106), .A2(gray_img[1408]), .B1(gray_img[1664]), .B2(
        n22770), .O(n22114) );
  MOAI1S U27675 ( .A1(n22797), .A2(intadd_62_B_0_), .B1(n22863), .B2(
        gray_img[1808]), .O(n22113) );
  AN4B1S U27676 ( .I1(n22116), .I2(n22115), .I3(n22114), .B1(n22113), .O(
        n22138) );
  AOI22S U27677 ( .A1(n22796), .A2(gray_img[1680]), .B1(gray_img[1424]), .B2(
        n22664), .O(n22124) );
  ND2S U27678 ( .I1(n22630), .I2(gray_img[512]), .O(n22121) );
  AOI22S U27679 ( .A1(gray_img[16]), .A2(n22901), .B1(gray_img[1936]), .B2(
        n22679), .O(n22120) );
  ND2S U27680 ( .I1(n22812), .I2(gray_img[1920]), .O(n22119) );
  NR2 U27681 ( .I1(n22117), .I2(n22811), .O(n22118) );
  AN4B1S U27682 ( .I1(n22121), .I2(n22120), .I3(n22119), .B1(n22118), .O(
        n22123) );
  AOI22S U27683 ( .A1(n22566), .A2(gray_img[896]), .B1(gray_img[640]), .B2(
        n22909), .O(n22122) );
  ND3S U27684 ( .I1(n22124), .I2(n22123), .I3(n22122), .O(n22131) );
  INV1S U27685 ( .I(gray_img[0]), .O(n23432) );
  NR2 U27686 ( .I1(n23432), .I2(n22125), .O(n22130) );
  AOI22S U27687 ( .A1(n21090), .A2(gray_img[1176]), .B1(n21137), .B2(
        gray_img[24]), .O(n22128) );
  AOI22S U27688 ( .A1(n22847), .A2(gray_img[1416]), .B1(n22619), .B2(
        gray_img[400]), .O(n22127) );
  AOI22S U27689 ( .A1(n22695), .A2(gray_img[656]), .B1(gray_img[912]), .B2(
        n22894), .O(n22126) );
  ND3S U27690 ( .I1(n22128), .I2(n22127), .I3(n22126), .O(n22129) );
  NR3 U27691 ( .I1(n22131), .I2(n22130), .I3(n22129), .O(n22137) );
  AOI22S U27692 ( .A1(n15915), .A2(gray_img[528]), .B1(gray_img[784]), .B2(
        n22930), .O(n22136) );
  ND2S U27693 ( .I1(n22929), .I2(gray_img[1040]), .O(n22134) );
  AOI22S U27694 ( .A1(n22625), .A2(gray_img[256]), .B1(gray_img[768]), .B2(
        n22513), .O(n22133) );
  AOI22S U27695 ( .A1(n22610), .A2(gray_img[128]), .B1(gray_img[776]), .B2(
        n22724), .O(n22132) );
  ND3S U27696 ( .I1(n22134), .I2(n22133), .I3(n22132), .O(n22135) );
  AN4B1S U27697 ( .I1(n22138), .I2(n22137), .I3(n22136), .B1(n22135), .O(
        n22152) );
  AOI22S U27698 ( .A1(n21155), .A2(gray_img[1032]), .B1(gray_img[1544]), .B2(
        n22656), .O(n22143) );
  AOI22S U27699 ( .A1(n22935), .A2(gray_img[1048]), .B1(gray_img[1816]), .B2(
        n22787), .O(n22142) );
  AOI22S U27700 ( .A1(n22837), .A2(gray_img[264]), .B1(gray_img[136]), .B2(
        n22933), .O(n22141) );
  INV1S U27701 ( .I(gray_img[1792]), .O(n22139) );
  MOAI1S U27702 ( .A1(n22364), .A2(n22139), .B1(n22934), .B2(gray_img[1280]), 
        .O(n22140) );
  AN4B1S U27703 ( .I1(n22143), .I2(n22142), .I3(n22141), .B1(n22140), .O(
        n22151) );
  ND2S U27704 ( .I1(n22931), .I2(gray_img[1928]), .O(n22150) );
  AOI22S U27705 ( .A1(n22867), .A2(gray_img[792]), .B1(gray_img[152]), .B2(
        n21089), .O(n22145) );
  AOI22S U27706 ( .A1(n22846), .A2(gray_img[1288]), .B1(gray_img[1800]), .B2(
        n22937), .O(n22144) );
  OA112S U27707 ( .C1(n29064), .C2(n22750), .A1(n22145), .B1(n22144), .O(
        n22148) );
  AOI22S U27708 ( .A1(n21096), .A2(gray_img[1432]), .B1(gray_img[1560]), .B2(
        n22918), .O(n22147) );
  ND2S U27709 ( .I1(n22755), .I2(gray_img[1944]), .O(n22146) );
  AN4B1S U27710 ( .I1(n22152), .I2(n22151), .I3(n22150), .B1(n22149), .O(
        n22153) );
  AOI22S U27711 ( .A1(n21152), .A2(gray_img[632]), .B1(gray_img[1656]), .B2(
        n22918), .O(n22160) );
  AOI22S U27712 ( .A1(n22724), .A2(gray_img[872]), .B1(n15921), .B2(
        gray_img[1264]), .O(n22159) );
  AOI22S U27713 ( .A1(n22786), .A2(gray_img[1784]), .B1(gray_img[864]), .B2(
        n22513), .O(n22158) );
  MOAI1S U27714 ( .A1(n22156), .A2(n26161), .B1(n22795), .B2(gray_img[616]), 
        .O(n22157) );
  AN4B1S U27715 ( .I1(n22160), .I2(n22159), .I3(n22158), .B1(n22157), .O(
        n22213) );
  ND2S U27716 ( .I1(n22867), .I2(gray_img[888]), .O(n22166) );
  AOI22S U27717 ( .A1(gray_img[1272]), .A2(n21090), .B1(n22881), .B2(
        gray_img[504]), .O(n22165) );
  ND2S U27718 ( .I1(n22889), .I2(gray_img[1392]), .O(n22164) );
  AOI22S U27719 ( .A1(n22935), .A2(gray_img[1144]), .B1(gray_img[1640]), .B2(
        n22874), .O(n22162) );
  AOI22S U27720 ( .A1(n22785), .A2(gray_img[376]), .B1(gray_img[352]), .B2(
        n22625), .O(n22161) );
  ND2S U27721 ( .I1(n22162), .I2(n22161), .O(n22163) );
  AN4B1S U27722 ( .I1(n22166), .I2(n22165), .I3(n22164), .B1(n22163), .O(
        n22212) );
  ND2S U27723 ( .I1(n22929), .I2(gray_img[1136]), .O(n22173) );
  AOI22S U27724 ( .A1(n22837), .A2(gray_img[360]), .B1(gray_img[232]), .B2(
        n22933), .O(n22172) );
  AOI22S U27725 ( .A1(n22864), .A2(gray_img[1912]), .B1(gray_img[1376]), .B2(
        n22934), .O(n22171) );
  ND2S U27726 ( .I1(n22930), .I2(gray_img[880]), .O(n22169) );
  AOI22S U27727 ( .A1(n21097), .A2(gray_img[1632]), .B1(gray_img[1248]), .B2(
        n22838), .O(n22168) );
  AOI22S U27728 ( .A1(n22610), .A2(gray_img[224]), .B1(gray_img[488]), .B2(
        n22862), .O(n22167) );
  AN4B1S U27729 ( .I1(n22173), .I2(n22172), .I3(n22171), .B1(n22170), .O(
        n22181) );
  AOI22S U27730 ( .A1(n21155), .A2(gray_img[1128]), .B1(gray_img[1256]), .B2(
        n22936), .O(n22179) );
  AOI22S U27731 ( .A1(n22861), .A2(gray_img[1384]), .B1(gray_img[1768]), .B2(
        n22921), .O(n22178) );
  AOI22S U27732 ( .A1(n22938), .A2(gray_img[1888]), .B1(gray_img[1120]), .B2(
        n22703), .O(n22177) );
  INV1S U27733 ( .I(gray_img[1896]), .O(n22174) );
  MOAI1S U27734 ( .A1(n22175), .A2(n22174), .B1(n22369), .B2(gray_img[1512]), 
        .O(n22176) );
  AN4B1S U27735 ( .I1(n22179), .I2(n22178), .I3(n22177), .B1(n22176), .O(
        n22180) );
  OAI112HS U27736 ( .C1(intadd_5_B_0_), .C2(n22853), .A1(n22181), .B1(n22180), 
        .O(n22210) );
  AOI22S U27737 ( .A1(n22695), .A2(gray_img[752]), .B1(gray_img[1008]), .B2(
        n22894), .O(n22186) );
  AOI22S U27738 ( .A1(n22619), .A2(gray_img[496]), .B1(gray_img[1776]), .B2(
        n22896), .O(n22185) );
  ND2S U27739 ( .I1(n21137), .I2(gray_img[120]), .O(n22184) );
  MOAI1S U27740 ( .A1(n22601), .A2(n22182), .B1(n22664), .B2(gray_img[1520]), 
        .O(n22183) );
  AN4B1S U27741 ( .I1(n22186), .I2(n22185), .I3(n22184), .B1(n22183), .O(
        n22189) );
  AOI22S U27742 ( .A1(n21096), .A2(gray_img[1528]), .B1(gray_img[1400]), .B2(
        n21120), .O(n22188) );
  ND2S U27743 ( .I1(n22919), .I2(gray_img[2040]), .O(n22187) );
  ND3S U27744 ( .I1(n22189), .I2(n22188), .I3(n22187), .O(n22209) );
  AOI22S U27745 ( .A1(n15905), .A2(gray_img[368]), .B1(gray_img[624]), .B2(
        n15915), .O(n22195) );
  MOAI1S U27746 ( .A1(n22346), .A2(n22190), .B1(n22883), .B2(gray_img[760]), 
        .O(n22192) );
  INV1S U27747 ( .I(gray_img[1504]), .O(n27985) );
  MOAI1S U27748 ( .A1(n22718), .A2(n27985), .B1(n22770), .B2(gray_img[1760]), 
        .O(n22191) );
  NR2 U27749 ( .I1(n22192), .I2(n22191), .O(n22194) );
  ND2S U27750 ( .I1(n15918), .I2(gray_img[240]), .O(n22193) );
  ND3S U27751 ( .I1(n22195), .I2(n22194), .I3(n22193), .O(n22207) );
  AOI22S U27752 ( .A1(n22630), .A2(gray_img[608]), .B1(gray_img[480]), .B2(
        n22686), .O(n22202) );
  ND2S U27753 ( .I1(n22819), .I2(gray_img[1016]), .O(n22201) );
  ND2S U27754 ( .I1(n22900), .I2(gray_img[104]), .O(n22200) );
  ND2S U27755 ( .I1(n22812), .I2(gray_img[2016]), .O(n22198) );
  AOI22S U27756 ( .A1(gray_img[248]), .A2(n21089), .B1(gray_img[2032]), .B2(
        n22679), .O(n22197) );
  ND2S U27757 ( .I1(gray_img[112]), .I2(n22901), .O(n22196) );
  AN4B1S U27758 ( .I1(n22202), .I2(n22201), .I3(n22200), .B1(n22199), .O(
        n22205) );
  AOI22S U27759 ( .A1(n22566), .A2(gray_img[992]), .B1(gray_img[744]), .B2(
        n22888), .O(n22204) );
  ND2S U27760 ( .I1(n22863), .I2(gray_img[1904]), .O(n22203) );
  ND3S U27761 ( .I1(n22205), .I2(n22204), .I3(n22203), .O(n22206) );
  AO112S U27762 ( .C1(gray_img[96]), .C2(n22893), .A1(n22207), .B1(n22206), 
        .O(n22208) );
  NR3 U27763 ( .I1(n22210), .I2(n22209), .I3(n22208), .O(n22211) );
  ND3S U27764 ( .I1(n22213), .I2(n22212), .I3(n22211), .O(n22214) );
  AOI22S U27765 ( .A1(n22784), .A2(n22215), .B1(n22959), .B2(n22214), .O(
        n22216) );
  INV1S U27766 ( .I(gray_img[1130]), .O(n28045) );
  MOAI1S U27767 ( .A1(n22848), .A2(n28045), .B1(n22864), .B2(gray_img[1914]), 
        .O(n22224) );
  INV1S U27768 ( .I(gray_img[1642]), .O(n25782) );
  MOAI1S U27769 ( .A1(n22218), .A2(n25782), .B1(n22861), .B2(gray_img[1386]), 
        .O(n22223) );
  ND2S U27770 ( .I1(n21152), .I2(gray_img[634]), .O(n22221) );
  AOI22S U27771 ( .A1(gray_img[370]), .A2(n15905), .B1(n22911), .B2(
        gray_img[994]), .O(n22220) );
  ND2S U27772 ( .I1(n22664), .I2(gray_img[1522]), .O(n22219) );
  ND3S U27773 ( .I1(n22221), .I2(n22220), .I3(n22219), .O(n22222) );
  NR3 U27774 ( .I1(n22224), .I2(n22223), .I3(n22222), .O(n22272) );
  ND2S U27775 ( .I1(n15915), .I2(gray_img[626]), .O(n22230) );
  AOI22S U27776 ( .A1(n22921), .A2(gray_img[1770]), .B1(n22827), .B2(
        gray_img[1650]), .O(n22229) );
  ND2S U27777 ( .I1(n21090), .I2(gray_img[1274]), .O(n22228) );
  AOI22S U27778 ( .A1(n22770), .A2(gray_img[1762]), .B1(n22703), .B2(
        gray_img[1122]), .O(n22226) );
  AOI22S U27779 ( .A1(gray_img[882]), .A2(n22930), .B1(n22810), .B2(
        gray_img[738]), .O(n22225) );
  ND2S U27780 ( .I1(n22226), .I2(n22225), .O(n22227) );
  AN4B1S U27781 ( .I1(n22230), .I2(n22229), .I3(n22228), .B1(n22227), .O(
        n22271) );
  ND2S U27782 ( .I1(n22893), .I2(gray_img[98]), .O(n22233) );
  AOI22S U27783 ( .A1(n22847), .A2(gray_img[1514]), .B1(n22619), .B2(
        gray_img[498]), .O(n22232) );
  AOI22S U27784 ( .A1(n22695), .A2(gray_img[754]), .B1(gray_img[1010]), .B2(
        n22894), .O(n22231) );
  ND3S U27785 ( .I1(n22233), .I2(n22232), .I3(n22231), .O(n22254) );
  AOI22S U27786 ( .A1(n22802), .A2(gray_img[1002]), .B1(gray_img[618]), .B2(
        n22795), .O(n22237) );
  ND2S U27787 ( .I1(n22863), .I2(gray_img[1906]), .O(n22236) );
  AOI22S U27788 ( .A1(n22657), .A2(gray_img[746]), .B1(gray_img[1786]), .B2(
        n22505), .O(n22235) );
  INV1S U27789 ( .I(gray_img[1394]), .O(n27907) );
  NR2 U27790 ( .I1(n27907), .I2(n22797), .O(n22234) );
  AN4B1S U27791 ( .I1(n22237), .I2(n22236), .I3(n22235), .B1(n22234), .O(
        n22246) );
  AOI22S U27792 ( .A1(n22630), .A2(gray_img[610]), .B1(gray_img[482]), .B2(
        n22686), .O(n22243) );
  ND2S U27793 ( .I1(n22819), .I2(gray_img[1018]), .O(n22242) );
  ND2S U27794 ( .I1(n22900), .I2(gray_img[106]), .O(n22241) );
  AOI22S U27795 ( .A1(gray_img[1530]), .A2(n21096), .B1(gray_img[2034]), .B2(
        n22679), .O(n22239) );
  ND2S U27796 ( .I1(gray_img[114]), .I2(n22901), .O(n22238) );
  OAI112HS U27797 ( .C1(n22904), .C2(n25838), .A1(n22239), .B1(n22238), .O(
        n22240) );
  AN4B1S U27798 ( .I1(n22243), .I2(n22242), .I3(n22241), .B1(n22240), .O(
        n22245) );
  AOI22S U27799 ( .A1(n22796), .A2(gray_img[1778]), .B1(gray_img[1266]), .B2(
        n15921), .O(n22244) );
  INV1S U27800 ( .I(gray_img[2042]), .O(n25947) );
  AOI22S U27801 ( .A1(n21089), .A2(gray_img[250]), .B1(gray_img[1658]), .B2(
        n22918), .O(n22248) );
  AOI22S U27802 ( .A1(n22727), .A2(gray_img[1898]), .B1(gray_img[1258]), .B2(
        n22936), .O(n22247) );
  AOI22S U27803 ( .A1(n21120), .A2(gray_img[1402]), .B1(n21137), .B2(
        gray_img[122]), .O(n22249) );
  OAI112HS U27804 ( .C1(n25947), .C2(n22251), .A1(n22250), .B1(n22249), .O(
        n22252) );
  NR3 U27805 ( .I1(n22254), .I2(n22253), .I3(n22252), .O(n22269) );
  AOI22S U27806 ( .A1(n22883), .A2(gray_img[762]), .B1(gray_img[378]), .B2(
        n22735), .O(n22258) );
  AOI22S U27807 ( .A1(n22625), .A2(gray_img[354]), .B1(gray_img[226]), .B2(
        n22610), .O(n22257) );
  AOI22S U27808 ( .A1(n22736), .A2(gray_img[506]), .B1(gray_img[1506]), .B2(
        n21106), .O(n22256) );
  INV1S U27809 ( .I(gray_img[1634]), .O(n25794) );
  MOAI1S U27810 ( .A1(n22670), .A2(n25794), .B1(n22872), .B2(gray_img[1250]), 
        .O(n22255) );
  AN4B1S U27811 ( .I1(n22258), .I2(n22257), .I3(n22256), .B1(n22255), .O(
        n22268) );
  ND2S U27812 ( .I1(n22663), .I2(gray_img[1138]), .O(n22262) );
  AOI22S U27813 ( .A1(n22836), .A2(gray_img[234]), .B1(gray_img[1146]), .B2(
        n22935), .O(n22261) );
  AOI22S U27814 ( .A1(n22938), .A2(gray_img[1890]), .B1(gray_img[1378]), .B2(
        n22934), .O(n22260) );
  NR2 U27815 ( .I1(n25850), .I2(n22853), .O(n22259) );
  AN4B1S U27816 ( .I1(n22262), .I2(n22261), .I3(n22260), .B1(n22259), .O(
        n22267) );
  ND2S U27817 ( .I1(n15918), .I2(gray_img[242]), .O(n22265) );
  AOI22S U27818 ( .A1(n22513), .A2(gray_img[866]), .B1(gray_img[362]), .B2(
        n22837), .O(n22264) );
  AOI22S U27819 ( .A1(n22724), .A2(gray_img[874]), .B1(gray_img[490]), .B2(
        n22862), .O(n22263) );
  ND3S U27820 ( .I1(n22265), .I2(n22264), .I3(n22263), .O(n22266) );
  AN4B1S U27821 ( .I1(n22269), .I2(n22268), .I3(n22267), .B1(n22266), .O(
        n22270) );
  ND2S U27822 ( .I1(n15918), .I2(gray_img[210]), .O(n22278) );
  AOI22S U27823 ( .A1(n22935), .A2(gray_img[1114]), .B1(gray_img[1738]), .B2(
        n22921), .O(n22277) );
  ND2S U27824 ( .I1(n21096), .I2(gray_img[1498]), .O(n22276) );
  AOI22S U27825 ( .A1(n22881), .A2(gray_img[474]), .B1(gray_img[842]), .B2(
        n22932), .O(n22274) );
  AOI22S U27826 ( .A1(gray_img[858]), .A2(n22813), .B1(n22786), .B2(
        gray_img[1754]), .O(n22273) );
  ND2S U27827 ( .I1(n22274), .I2(n22273), .O(n22275) );
  AN4B1S U27828 ( .I1(n22278), .I2(n22277), .I3(n22276), .B1(n22275), .O(
        n22324) );
  AOI22S U27829 ( .A1(n22695), .A2(gray_img[722]), .B1(gray_img[1234]), .B2(
        n15921), .O(n22282) );
  AOI22S U27830 ( .A1(gray_img[594]), .A2(n15915), .B1(n22873), .B2(
        gray_img[986]), .O(n22281) );
  AOI22S U27831 ( .A1(n22872), .A2(gray_img[1218]), .B1(gray_img[330]), .B2(
        n22837), .O(n22280) );
  INV1S U27832 ( .I(gray_img[1098]), .O(n28483) );
  MOAI1S U27833 ( .A1(n28483), .A2(n22848), .B1(n22828), .B2(gray_img[978]), 
        .O(n22279) );
  AN4B1S U27834 ( .I1(n22282), .I2(n22281), .I3(n22280), .B1(n22279), .O(
        n22323) );
  ND2S U27835 ( .I1(n22893), .I2(gray_img[66]), .O(n22285) );
  AOI22S U27836 ( .A1(n22874), .A2(gray_img[1610]), .B1(n22619), .B2(
        gray_img[466]), .O(n22284) );
  AOI22S U27837 ( .A1(n22796), .A2(gray_img[1746]), .B1(gray_img[1490]), .B2(
        n22664), .O(n22283) );
  ND3S U27838 ( .I1(n22285), .I2(n22284), .I3(n22283), .O(n22301) );
  ND2S U27839 ( .I1(n22827), .I2(gray_img[1618]), .O(n22291) );
  ND2S U27840 ( .I1(n22909), .I2(gray_img[706]), .O(n22290) );
  ND2S U27841 ( .I1(n22812), .I2(gray_img[1986]), .O(n22289) );
  INV1S U27842 ( .I(gray_img[74]), .O(n23591) );
  AOI22S U27843 ( .A1(gray_img[2002]), .A2(n22679), .B1(gray_img[1370]), .B2(
        n21120), .O(n22287) );
  AOI22S U27844 ( .A1(gray_img[1626]), .A2(n22918), .B1(gray_img[82]), .B2(
        n22901), .O(n22286) );
  OAI112HS U27845 ( .C1(n22811), .C2(n23591), .A1(n22287), .B1(n22286), .O(
        n22288) );
  AN4B1S U27846 ( .I1(n22291), .I2(n22290), .I3(n22289), .B1(n22288), .O(
        n22294) );
  AOI22S U27847 ( .A1(n22566), .A2(gray_img[962]), .B1(gray_img[450]), .B2(
        n22686), .O(n22293) );
  AOI22S U27848 ( .A1(n22630), .A2(gray_img[578]), .B1(gray_img[970]), .B2(
        n22910), .O(n22292) );
  ND3S U27849 ( .I1(n22294), .I2(n22293), .I3(n22292), .O(n22300) );
  INV1S U27850 ( .I(gray_img[1362]), .O(n28374) );
  AOI22S U27851 ( .A1(n22657), .A2(gray_img[714]), .B1(gray_img[586]), .B2(
        n22795), .O(n22295) );
  AOI22S U27852 ( .A1(n22883), .A2(gray_img[730]), .B1(gray_img[346]), .B2(
        n22735), .O(n22297) );
  ND2S U27853 ( .I1(n22863), .I2(gray_img[1874]), .O(n22296) );
  ND3S U27854 ( .I1(n22298), .I2(n22297), .I3(n22296), .O(n22299) );
  NR3 U27855 ( .I1(n22301), .I2(n22300), .I3(n22299), .O(n22308) );
  AOI22S U27856 ( .A1(n21090), .A2(gray_img[1242]), .B1(n21137), .B2(
        gray_img[90]), .O(n22307) );
  ND2S U27857 ( .I1(n22755), .I2(gray_img[2010]), .O(n22306) );
  AOI22S U27858 ( .A1(n21152), .A2(gray_img[602]), .B1(gray_img[218]), .B2(
        n21089), .O(n22304) );
  AOI22S U27859 ( .A1(n22847), .A2(gray_img[1482]), .B1(gray_img[1226]), .B2(
        n22936), .O(n22303) );
  AOI22S U27860 ( .A1(n22846), .A2(gray_img[1354]), .B1(gray_img[1866]), .B2(
        n22727), .O(n22302) );
  ND3S U27861 ( .I1(n22304), .I2(n22303), .I3(n22302), .O(n22305) );
  AN4B1S U27862 ( .I1(n22308), .I2(n22307), .I3(n22306), .B1(n22305), .O(
        n22321) );
  AOI22S U27863 ( .A1(n21106), .A2(gray_img[1474]), .B1(gray_img[1602]), .B2(
        n21097), .O(n22314) );
  AOI22S U27864 ( .A1(n22770), .A2(gray_img[1730]), .B1(gray_img[834]), .B2(
        n22513), .O(n22313) );
  ND2S U27865 ( .I1(n15905), .I2(gray_img[338]), .O(n22312) );
  AOI22S U27866 ( .A1(n22625), .A2(gray_img[322]), .B1(gray_img[194]), .B2(
        n22610), .O(n22310) );
  AOI22S U27867 ( .A1(n22933), .A2(gray_img[202]), .B1(gray_img[458]), .B2(
        n22762), .O(n22309) );
  OAI112HS U27868 ( .C1(n22841), .C2(intadd_97_B_1_), .A1(n22310), .B1(n22309), 
        .O(n22311) );
  AN4B1S U27869 ( .I1(n22314), .I2(n22313), .I3(n22312), .B1(n22311), .O(
        n22320) );
  ND2S U27870 ( .I1(n22931), .I2(gray_img[1994]), .O(n22319) );
  ND2S U27871 ( .I1(n22663), .I2(gray_img[1106]), .O(n22317) );
  AOI22S U27872 ( .A1(n22864), .A2(gray_img[1882]), .B1(gray_img[1090]), .B2(
        n22703), .O(n22316) );
  AOI22S U27873 ( .A1(n22938), .A2(gray_img[1858]), .B1(gray_img[1346]), .B2(
        n22934), .O(n22315) );
  ND3S U27874 ( .I1(n22317), .I2(n22316), .I3(n22315), .O(n22318) );
  AN4B1S U27875 ( .I1(n22321), .I2(n22320), .I3(n22319), .B1(n22318), .O(
        n22322) );
  AOI22S U27876 ( .A1(n22959), .A2(n22326), .B1(n22782), .B2(n22325), .O(
        n22435) );
  AOI22S U27877 ( .A1(n22770), .A2(gray_img[1666]), .B1(n15921), .B2(
        gray_img[1170]), .O(n22330) );
  AOI22S U27878 ( .A1(gray_img[1434]), .A2(n21096), .B1(n22566), .B2(
        gray_img[898]), .O(n22329) );
  AOI22S U27879 ( .A1(n22810), .A2(gray_img[642]), .B1(gray_img[666]), .B2(
        n22883), .O(n22328) );
  INV1S U27880 ( .I(gray_img[1682]), .O(n26548) );
  MOAI1S U27881 ( .A1(n22540), .A2(n26548), .B1(n22827), .B2(gray_img[1554]), 
        .O(n22327) );
  AN4B1S U27882 ( .I1(n22330), .I2(n22329), .I3(n22328), .B1(n22327), .O(
        n22379) );
  MOAI1S U27883 ( .A1(n22392), .A2(n26629), .B1(n22935), .B2(gray_img[1050]), 
        .O(n22335) );
  INV1S U27884 ( .I(gray_img[1674]), .O(n26577) );
  MOAI1S U27885 ( .A1(n22487), .A2(n26577), .B1(n22727), .B2(gray_img[1802]), 
        .O(n22334) );
  ND2S U27886 ( .I1(n21120), .I2(gray_img[1306]), .O(n22332) );
  AOI22S U27887 ( .A1(n22686), .A2(gray_img[386]), .B1(gray_img[650]), .B2(
        n22657), .O(n22331) );
  OAI112HS U27888 ( .C1(n22848), .C2(intadd_89_B_1_), .A1(n22332), .B1(n22331), 
        .O(n22333) );
  NR3 U27889 ( .I1(n22335), .I2(n22334), .I3(n22333), .O(n22378) );
  AOI22S U27890 ( .A1(n22785), .A2(gray_img[282]), .B1(gray_img[410]), .B2(
        n22881), .O(n22339) );
  ND2S U27891 ( .I1(n22863), .I2(gray_img[1810]), .O(n22338) );
  AOI22S U27892 ( .A1(n22795), .A2(gray_img[522]), .B1(gray_img[1690]), .B2(
        n22505), .O(n22337) );
  INV1S U27893 ( .I(gray_img[1410]), .O(n29646) );
  MOAI1S U27894 ( .A1(n22718), .A2(n29646), .B1(n21097), .B2(gray_img[1538]), 
        .O(n22336) );
  AN4B1S U27895 ( .I1(n22339), .I2(n22338), .I3(n22337), .B1(n22336), .O(
        n22352) );
  AOI22S U27896 ( .A1(n15918), .A2(gray_img[146]), .B1(gray_img[530]), .B2(
        n15915), .O(n22351) );
  AOI22S U27897 ( .A1(n15905), .A2(gray_img[274]), .B1(gray_img[786]), .B2(
        n22930), .O(n22350) );
  INV1S U27898 ( .I(gray_img[922]), .O(n29276) );
  ND2S U27899 ( .I1(n22664), .I2(gray_img[1426]), .O(n22345) );
  ND2S U27900 ( .I1(n22812), .I2(gray_img[1922]), .O(n22343) );
  AOI22S U27901 ( .A1(gray_img[1938]), .A2(n22679), .B1(gray_img[154]), .B2(
        n21089), .O(n22342) );
  ND2S U27902 ( .I1(gray_img[18]), .I2(n22901), .O(n22341) );
  INV1S U27903 ( .I(gray_img[10]), .O(n23420) );
  NR2 U27904 ( .I1(n23420), .I2(n22811), .O(n22340) );
  AN4B1S U27905 ( .I1(n22343), .I2(n22342), .I3(n22341), .B1(n22340), .O(
        n22344) );
  OAI112HS U27906 ( .C1(n22682), .C2(n29276), .A1(n22345), .B1(n22344), .O(
        n22348) );
  MOAI1S U27907 ( .A1(n22346), .A2(n29606), .B1(n22630), .B2(gray_img[514]), 
        .O(n22347) );
  AO112S U27908 ( .C1(gray_img[1298]), .C2(n22889), .A1(n22348), .B1(n22347), 
        .O(n22349) );
  AN4B1S U27909 ( .I1(n22352), .I2(n22351), .I3(n22350), .B1(n22349), .O(
        n22359) );
  AOI22S U27910 ( .A1(n21090), .A2(gray_img[1178]), .B1(n21137), .B2(
        gray_img[26]), .O(n22358) );
  ND2S U27911 ( .I1(n22755), .I2(gray_img[1946]), .O(n22357) );
  ND2S U27912 ( .I1(n22893), .I2(gray_img[2]), .O(n22355) );
  AOI22S U27913 ( .A1(n22936), .A2(gray_img[1162]), .B1(n22619), .B2(
        gray_img[402]), .O(n22354) );
  AOI22S U27914 ( .A1(n22695), .A2(gray_img[658]), .B1(gray_img[914]), .B2(
        n22894), .O(n22353) );
  ND3S U27915 ( .I1(n22355), .I2(n22354), .I3(n22353), .O(n22356) );
  AN4B1S U27916 ( .I1(n22359), .I2(n22358), .I3(n22357), .B1(n22356), .O(
        n22376) );
  ND2S U27917 ( .I1(n22663), .I2(gray_img[1042]), .O(n22363) );
  AOI22S U27918 ( .A1(n22513), .A2(gray_img[770]), .B1(gray_img[130]), .B2(
        n22610), .O(n22362) );
  AOI22S U27919 ( .A1(n22625), .A2(gray_img[258]), .B1(gray_img[778]), .B2(
        n22724), .O(n22361) );
  NR2 U27920 ( .I1(n29402), .I2(n22853), .O(n22360) );
  AN4B1S U27921 ( .I1(n22363), .I2(n22362), .I3(n22361), .B1(n22360), .O(
        n22375) );
  AOI22S U27922 ( .A1(n22703), .A2(gray_img[1026]), .B1(gray_img[1546]), .B2(
        n22656), .O(n22368) );
  AOI22S U27923 ( .A1(n22837), .A2(gray_img[266]), .B1(gray_img[394]), .B2(
        n22862), .O(n22367) );
  AOI22S U27924 ( .A1(n22836), .A2(gray_img[138]), .B1(gray_img[1818]), .B2(
        n22787), .O(n22366) );
  INV1S U27925 ( .I(gray_img[1794]), .O(n29389) );
  MOAI1S U27926 ( .A1(n22364), .A2(n29389), .B1(n22934), .B2(gray_img[1282]), 
        .O(n22365) );
  AN4B1S U27927 ( .I1(n22368), .I2(n22367), .I3(n22366), .B1(n22365), .O(
        n22374) );
  AOI22S U27928 ( .A1(n22813), .A2(gray_img[794]), .B1(gray_img[1562]), .B2(
        n22918), .O(n22372) );
  AOI22S U27929 ( .A1(n22846), .A2(gray_img[1290]), .B1(gray_img[1418]), .B2(
        n22369), .O(n22371) );
  ND2S U27930 ( .I1(n21152), .I2(gray_img[538]), .O(n22370) );
  AN4B1S U27931 ( .I1(n22376), .I2(n22375), .I3(n22374), .B1(n22373), .O(
        n22377) );
  NR2 U27932 ( .I1(n22380), .I2(n22493), .O(n22386) );
  INV1S U27933 ( .I(gray_img[1714]), .O(n29211) );
  MOAI1S U27934 ( .A1(n22540), .A2(n29211), .B1(gray_img[1194]), .B2(n22936), 
        .O(n22385) );
  INV1S U27935 ( .I(gray_img[306]), .O(n26503) );
  AOI22S U27936 ( .A1(gray_img[1074]), .A2(n22929), .B1(n22887), .B2(
        gray_img[554]), .O(n22382) );
  AOI22S U27937 ( .A1(n22802), .A2(gray_img[938]), .B1(gray_img[802]), .B2(
        n22513), .O(n22381) );
  OAI112HS U27938 ( .C1(n22383), .C2(n26503), .A1(n22382), .B1(n22381), .O(
        n22384) );
  NR3 U27939 ( .I1(n22386), .I2(n22385), .I3(n22384), .O(n22431) );
  AOI22S U27940 ( .A1(n22813), .A2(gray_img[826]), .B1(gray_img[186]), .B2(
        n21089), .O(n22391) );
  AOI22S U27941 ( .A1(gray_img[818]), .A2(n22930), .B1(n22657), .B2(
        gray_img[682]), .O(n22390) );
  ND2S U27942 ( .I1(n15921), .I2(gray_img[1202]), .O(n22389) );
  INV1S U27943 ( .I(gray_img[1442]), .O(n28952) );
  MOAI1S U27944 ( .A1(n22718), .A2(n28952), .B1(n22864), .B2(gray_img[1850]), 
        .O(n22387) );
  AO12S U27945 ( .B1(gray_img[1330]), .B2(n22889), .A1(n22387), .O(n22388) );
  AN4B1S U27946 ( .I1(n22391), .I2(n22390), .I3(n22389), .B1(n22388), .O(
        n22430) );
  AOI22S U27947 ( .A1(n22785), .A2(gray_img[314]), .B1(gray_img[442]), .B2(
        n22736), .O(n22396) );
  AOI22S U27948 ( .A1(n22770), .A2(gray_img[1698]), .B1(gray_img[290]), .B2(
        n22625), .O(n22395) );
  AOI22S U27949 ( .A1(n22786), .A2(gray_img[1722]), .B1(gray_img[698]), .B2(
        n22883), .O(n22394) );
  MOAI1S U27950 ( .A1(n22392), .A2(n23010), .B1(n21097), .B2(gray_img[1570]), 
        .O(n22393) );
  AN4B1S U27951 ( .I1(n22396), .I2(n22395), .I3(n22394), .B1(n22393), .O(
        n22408) );
  AOI22S U27952 ( .A1(n22566), .A2(gray_img[930]), .B1(gray_img[418]), .B2(
        n22686), .O(n22407) );
  ND2S U27953 ( .I1(n22863), .I2(gray_img[1842]), .O(n22406) );
  INV1S U27954 ( .I(gray_img[954]), .O(n26113) );
  AOI22S U27955 ( .A1(n22630), .A2(gray_img[546]), .B1(gray_img[674]), .B2(
        n22909), .O(n22404) );
  AOI22S U27956 ( .A1(gray_img[50]), .A2(n22901), .B1(gray_img[1338]), .B2(
        n21120), .O(n22399) );
  AOI22S U27957 ( .A1(gray_img[1210]), .A2(n21090), .B1(gray_img[1970]), .B2(
        n22679), .O(n22398) );
  ND2S U27958 ( .I1(gray_img[1594]), .I2(n22694), .O(n22397) );
  ND3S U27959 ( .I1(n22399), .I2(n22398), .I3(n22397), .O(n22402) );
  INV1S U27960 ( .I(gray_img[42]), .O(n26958) );
  NR2 U27961 ( .I1(n26958), .I2(n22811), .O(n22401) );
  NR2 U27962 ( .I1(n26658), .I2(n22904), .O(n22400) );
  NR3 U27963 ( .I1(n22402), .I2(n22401), .I3(n22400), .O(n22403) );
  OAI112HS U27964 ( .C1(n22682), .C2(n26113), .A1(n22404), .B1(n22403), .O(
        n22405) );
  AN4B1S U27965 ( .I1(n22408), .I2(n22407), .I3(n22406), .B1(n22405), .O(
        n22428) );
  AOI22S U27966 ( .A1(n15918), .A2(gray_img[178]), .B1(gray_img[562]), .B2(
        n15915), .O(n22427) );
  AOI22S U27967 ( .A1(n22938), .A2(gray_img[1826]), .B1(gray_img[1314]), .B2(
        n22934), .O(n22412) );
  AOI22S U27968 ( .A1(n22724), .A2(gray_img[810]), .B1(gray_img[1082]), .B2(
        n22935), .O(n22411) );
  AOI22S U27969 ( .A1(n22610), .A2(gray_img[162]), .B1(gray_img[426]), .B2(
        n22862), .O(n22410) );
  INV1S U27970 ( .I(gray_img[298]), .O(n27277) );
  MOAI1S U27971 ( .A1(n22865), .A2(n27277), .B1(n22836), .B2(gray_img[170]), 
        .O(n22409) );
  AN4B1S U27972 ( .I1(n22412), .I2(n22411), .I3(n22410), .B1(n22409), .O(
        n22426) );
  AOI22S U27973 ( .A1(n22619), .A2(gray_img[434]), .B1(gray_img[690]), .B2(
        n22920), .O(n22418) );
  AOI22S U27974 ( .A1(n22664), .A2(gray_img[1458]), .B1(gray_img[1586]), .B2(
        n15919), .O(n22417) );
  ND2S U27975 ( .I1(n22893), .I2(gray_img[34]), .O(n22416) );
  INV1S U27976 ( .I(gray_img[58]), .O(n27711) );
  ND2S U27977 ( .I1(n22919), .I2(gray_img[1978]), .O(n22414) );
  AOI22S U27978 ( .A1(n22847), .A2(gray_img[1450]), .B1(n22828), .B2(
        gray_img[946]), .O(n22413) );
  OAI112HS U27979 ( .C1(n22924), .C2(n27711), .A1(n22414), .B1(n22413), .O(
        n22415) );
  AN4B1S U27980 ( .I1(n22418), .I2(n22417), .I3(n22416), .B1(n22415), .O(
        n22424) );
  AOI22S U27981 ( .A1(n21155), .A2(gray_img[1066]), .B1(gray_img[1834]), .B2(
        n22937), .O(n22422) );
  AOI22S U27982 ( .A1(n22861), .A2(gray_img[1322]), .B1(gray_img[1706]), .B2(
        n22921), .O(n22421) );
  AOI22S U27983 ( .A1(n22703), .A2(gray_img[1058]), .B1(gray_img[1578]), .B2(
        n22656), .O(n22420) );
  INV1S U27984 ( .I(gray_img[570]), .O(n28145) );
  NR2 U27985 ( .I1(n28145), .I2(n22750), .O(n22419) );
  AN4B1S U27986 ( .I1(n22422), .I2(n22421), .I3(n22420), .B1(n22419), .O(
        n22423) );
  OAI112HS U27987 ( .C1(n26671), .C2(n22853), .A1(n22424), .B1(n22423), .O(
        n22425) );
  AN4B1S U27988 ( .I1(n22428), .I2(n22427), .I3(n22426), .B1(n22425), .O(
        n22429) );
  ND3S U27989 ( .I1(n22431), .I2(n22430), .I3(n22429), .O(n22432) );
  AOI22S U27990 ( .A1(n22784), .A2(n22433), .B1(n22957), .B2(n22432), .O(
        n22434) );
  AOI22S U27991 ( .A1(n22724), .A2(gray_img[777]), .B1(n22664), .B2(
        gray_img[1425]), .O(n22439) );
  AOI22S U27992 ( .A1(gray_img[1177]), .A2(n21090), .B1(n22911), .B2(
        gray_img[897]), .O(n22438) );
  AOI22S U27993 ( .A1(n22810), .A2(gray_img[641]), .B1(gray_img[521]), .B2(
        n22795), .O(n22437) );
  MOAI1S U27994 ( .A1(n22718), .A2(intadd_66_CI), .B1(n22910), .B2(
        gray_img[905]), .O(n22436) );
  AN4B1S U27995 ( .I1(n22439), .I2(n22438), .I3(n22437), .B1(n22436), .O(
        n22484) );
  AOI22S U27996 ( .A1(n22867), .A2(gray_img[793]), .B1(gray_img[1433]), .B2(
        n21096), .O(n22443) );
  AOI22S U27997 ( .A1(n22938), .A2(gray_img[1793]), .B1(n22827), .B2(
        gray_img[1553]), .O(n22442) );
  AOI22S U27998 ( .A1(n22610), .A2(gray_img[129]), .B1(gray_img[137]), .B2(
        n22836), .O(n22441) );
  INV1S U27999 ( .I(gray_img[1689]), .O(n26530) );
  MOAI1S U28000 ( .A1(n22882), .A2(n26530), .B1(gray_img[1561]), .B2(n22694), 
        .O(n22440) );
  AN4B1S U28001 ( .I1(n22443), .I2(n22442), .I3(n22441), .B1(n22440), .O(
        n22483) );
  AOI22S U28002 ( .A1(n22785), .A2(gray_img[281]), .B1(gray_img[409]), .B2(
        n22736), .O(n22447) );
  ND2S U28003 ( .I1(n22863), .I2(gray_img[1809]), .O(n22446) );
  AOI22S U28004 ( .A1(n22657), .A2(gray_img[649]), .B1(gray_img[665]), .B2(
        n22883), .O(n22445) );
  MOAI1S U28005 ( .A1(n22670), .A2(n26588), .B1(n22872), .B2(gray_img[1153]), 
        .O(n22444) );
  AN4B1S U28006 ( .I1(n22447), .I2(n22446), .I3(n22445), .B1(n22444), .O(
        n22459) );
  AOI22S U28007 ( .A1(n15905), .A2(gray_img[273]), .B1(gray_img[785]), .B2(
        n22930), .O(n22458) );
  AOI22S U28008 ( .A1(n15918), .A2(gray_img[145]), .B1(gray_img[529]), .B2(
        n15915), .O(n22457) );
  INV1S U28009 ( .I(gray_img[921]), .O(n29274) );
  NR2 U28010 ( .I1(n29274), .I2(n22682), .O(n22452) );
  AOI22S U28011 ( .A1(gray_img[17]), .A2(n22901), .B1(gray_img[1937]), .B2(
        n22679), .O(n22449) );
  ND2S U28012 ( .I1(n22812), .I2(gray_img[1921]), .O(n22448) );
  OAI112HS U28013 ( .C1(n22811), .C2(n23418), .A1(n22449), .B1(n22448), .O(
        n22451) );
  NR2 U28014 ( .I1(intadd_50_CI), .I2(n22540), .O(n22450) );
  NR3 U28015 ( .I1(n22452), .I2(n22451), .I3(n22450), .O(n22455) );
  AOI22S U28016 ( .A1(n22630), .A2(gray_img[513]), .B1(gray_img[385]), .B2(
        n22686), .O(n22454) );
  ND2S U28017 ( .I1(n22889), .I2(gray_img[1297]), .O(n22453) );
  ND3S U28018 ( .I1(n22455), .I2(n22454), .I3(n22453), .O(n22456) );
  AN4B1S U28019 ( .I1(n22459), .I2(n22458), .I3(n22457), .B1(n22456), .O(
        n22466) );
  AOI22S U28020 ( .A1(n21120), .A2(gray_img[1305]), .B1(n21137), .B2(
        gray_img[25]), .O(n22465) );
  ND2S U28021 ( .I1(n22755), .I2(gray_img[1945]), .O(n22464) );
  ND2S U28022 ( .I1(n22893), .I2(gray_img[1]), .O(n22462) );
  AOI22S U28023 ( .A1(n22920), .A2(gray_img[657]), .B1(gray_img[913]), .B2(
        n22894), .O(n22461) );
  AOI22S U28024 ( .A1(n22619), .A2(gray_img[401]), .B1(gray_img[1169]), .B2(
        n15921), .O(n22460) );
  ND3S U28025 ( .I1(n22462), .I2(n22461), .I3(n22460), .O(n22463) );
  AN4B1S U28026 ( .I1(n22466), .I2(n22465), .I3(n22464), .B1(n22463), .O(
        n22481) );
  ND2S U28027 ( .I1(n22663), .I2(gray_img[1041]), .O(n22470) );
  AOI22S U28028 ( .A1(n22770), .A2(gray_img[1665]), .B1(gray_img[769]), .B2(
        n22513), .O(n22469) );
  AOI22S U28029 ( .A1(n22625), .A2(gray_img[257]), .B1(gray_img[265]), .B2(
        n22837), .O(n22468) );
  INV1S U28030 ( .I(gray_img[1929]), .O(n29400) );
  NR2 U28031 ( .I1(n29400), .I2(n22853), .O(n22467) );
  AN4B1S U28032 ( .I1(n22470), .I2(n22469), .I3(n22468), .B1(n22467), .O(
        n22480) );
  AOI22S U28033 ( .A1(n22934), .A2(gray_img[1281]), .B1(gray_img[1289]), .B2(
        n22861), .O(n22474) );
  AOI22S U28034 ( .A1(n22935), .A2(gray_img[1049]), .B1(gray_img[1025]), .B2(
        n22703), .O(n22473) );
  AOI22S U28035 ( .A1(n22762), .A2(gray_img[393]), .B1(gray_img[1817]), .B2(
        n22864), .O(n22472) );
  INV1S U28036 ( .I(gray_img[1673]), .O(n26575) );
  MOAI1S U28037 ( .A1(n22487), .A2(n26575), .B1(n22656), .B2(gray_img[1545]), 
        .O(n22471) );
  AN4B1S U28038 ( .I1(n22474), .I2(n22473), .I3(n22472), .B1(n22471), .O(
        n22479) );
  AOI22S U28039 ( .A1(n21152), .A2(gray_img[537]), .B1(gray_img[153]), .B2(
        n21089), .O(n22477) );
  AOI22S U28040 ( .A1(n22847), .A2(gray_img[1417]), .B1(gray_img[1161]), .B2(
        n22936), .O(n22476) );
  AOI22S U28041 ( .A1(n21155), .A2(gray_img[1033]), .B1(gray_img[1801]), .B2(
        n22937), .O(n22475) );
  ND3S U28042 ( .I1(n22477), .I2(n22476), .I3(n22475), .O(n22478) );
  AN4B1S U28043 ( .I1(n22481), .I2(n22480), .I3(n22479), .B1(n22478), .O(
        n22482) );
  AOI22S U28044 ( .A1(n22933), .A2(gray_img[169]), .B1(gray_img[1057]), .B2(
        n22703), .O(n22490) );
  ND2S U28045 ( .I1(n22867), .I2(gray_img[825]), .O(n22486) );
  AOI22S U28046 ( .A1(n22810), .A2(gray_img[673]), .B1(gray_img[697]), .B2(
        n22883), .O(n22485) );
  OAI112HS U28047 ( .C1(n22487), .C2(intadd_47_CI), .A1(n22486), .B1(n22485), 
        .O(n22489) );
  MOAI1S U28048 ( .A1(n22884), .A2(intadd_13_CI), .B1(n22610), .B2(
        gray_img[161]), .O(n22488) );
  AN3B2S U28049 ( .I1(n22490), .B1(n22489), .B2(n22488), .O(n22537) );
  AOI22S U28050 ( .A1(n22864), .A2(gray_img[1849]), .B1(gray_img[1825]), .B2(
        n22794), .O(n22496) );
  AOI22S U28051 ( .A1(n22686), .A2(gray_img[417]), .B1(gray_img[441]), .B2(
        n22881), .O(n22492) );
  ND2S U28052 ( .I1(n22656), .I2(gray_img[1577]), .O(n22491) );
  OAI112HS U28053 ( .C1(n22493), .C2(intadd_134_CI), .A1(n22492), .B1(n22491), 
        .O(n22495) );
  MOAI1S U28054 ( .A1(n22718), .A2(intadd_60_CI), .B1(n22932), .B2(
        gray_img[809]), .O(n22494) );
  AN3B2S U28055 ( .I1(n22496), .B1(n22495), .B2(n22494), .O(n22536) );
  AOI22S U28056 ( .A1(n15905), .A2(gray_img[305]), .B1(gray_img[817]), .B2(
        n22930), .O(n22512) );
  AOI22S U28057 ( .A1(n15918), .A2(gray_img[177]), .B1(gray_img[561]), .B2(
        n15915), .O(n22511) );
  AOI22S U28058 ( .A1(n22657), .A2(gray_img[681]), .B1(gray_img[553]), .B2(
        n22795), .O(n22504) );
  AOI22S U28059 ( .A1(n22630), .A2(gray_img[545]), .B1(gray_img[929]), .B2(
        n22911), .O(n22503) );
  ND2S U28060 ( .I1(n15919), .I2(gray_img[1585]), .O(n22502) );
  ND2S U28061 ( .I1(n22819), .I2(gray_img[953]), .O(n22500) );
  ND2S U28062 ( .I1(n22812), .I2(gray_img[1953]), .O(n22498) );
  AOI22S U28063 ( .A1(gray_img[49]), .A2(n22901), .B1(gray_img[1969]), .B2(
        n22679), .O(n22497) );
  OA112S U28064 ( .C1(n22750), .C2(intadd_189_A_0_), .A1(n22498), .B1(n22497), 
        .O(n22499) );
  OAI112HS U28065 ( .C1(n22811), .C2(intadd_22_CI), .A1(n22500), .B1(n22499), 
        .O(n22501) );
  AN4B1S U28066 ( .I1(n22504), .I2(n22503), .I3(n22502), .B1(n22501), .O(
        n22510) );
  AOI22S U28067 ( .A1(n22863), .A2(gray_img[1841]), .B1(gray_img[1329]), .B2(
        n22889), .O(n22508) );
  AOI22S U28068 ( .A1(n22802), .A2(gray_img[937]), .B1(gray_img[1721]), .B2(
        n22505), .O(n22507) );
  AOI22S U28069 ( .A1(n21097), .A2(gray_img[1569]), .B1(gray_img[1185]), .B2(
        n22838), .O(n22506) );
  ND3S U28070 ( .I1(n22508), .I2(n22507), .I3(n22506), .O(n22509) );
  AN4B1S U28071 ( .I1(n22512), .I2(n22511), .I3(n22510), .B1(n22509), .O(
        n22534) );
  ND2S U28072 ( .I1(n22663), .I2(gray_img[1073]), .O(n22517) );
  AOI22S U28073 ( .A1(n22770), .A2(gray_img[1697]), .B1(gray_img[801]), .B2(
        n22513), .O(n22516) );
  AOI22S U28074 ( .A1(n22625), .A2(gray_img[289]), .B1(gray_img[297]), .B2(
        n22837), .O(n22515) );
  NR2 U28075 ( .I1(n26669), .I2(n22853), .O(n22514) );
  AN4B1S U28076 ( .I1(n22517), .I2(n22516), .I3(n22515), .B1(n22514), .O(
        n22533) );
  AOI22S U28077 ( .A1(n22828), .A2(gray_img[945]), .B1(gray_img[1201]), .B2(
        n15921), .O(n22523) );
  AOI22S U28078 ( .A1(n22796), .A2(gray_img[1713]), .B1(gray_img[1457]), .B2(
        n22664), .O(n22522) );
  ND2S U28079 ( .I1(n22893), .I2(gray_img[33]), .O(n22521) );
  ND2S U28080 ( .I1(n22755), .I2(gray_img[1977]), .O(n22519) );
  AOI22S U28081 ( .A1(n22619), .A2(gray_img[433]), .B1(gray_img[689]), .B2(
        n22920), .O(n22518) );
  OAI112HS U28082 ( .C1(n22924), .C2(n27709), .A1(n22519), .B1(n22518), .O(
        n22520) );
  AN4B1S U28083 ( .I1(n22523), .I2(n22522), .I3(n22521), .B1(n22520), .O(
        n22532) );
  AOI22S U28084 ( .A1(n22937), .A2(gray_img[1833]), .B1(gray_img[1193]), .B2(
        n22936), .O(n22527) );
  AOI22S U28085 ( .A1(n22934), .A2(gray_img[1313]), .B1(gray_img[1321]), .B2(
        n22846), .O(n22526) );
  AOI22S U28086 ( .A1(n22862), .A2(gray_img[425]), .B1(gray_img[1081]), .B2(
        n22935), .O(n22525) );
  MOAI1S U28087 ( .A1(n22875), .A2(intadd_59_CI), .B1(n21155), .B2(
        gray_img[1065]), .O(n22524) );
  AN4B1S U28088 ( .I1(n22527), .I2(n22526), .I3(n22525), .B1(n22524), .O(
        n22530) );
  AOI22S U28089 ( .A1(n21089), .A2(gray_img[185]), .B1(gray_img[1593]), .B2(
        n22918), .O(n22529) );
  AOI22S U28090 ( .A1(n21090), .A2(gray_img[1209]), .B1(gray_img[1337]), .B2(
        n21120), .O(n22528) );
  AN4B1S U28091 ( .I1(n22534), .I2(n22533), .I3(n22532), .B1(n22531), .O(
        n22535) );
  ND3S U28092 ( .I1(n22537), .I2(n22536), .I3(n22535), .O(n22538) );
  AOI22S U28093 ( .A1(n22784), .A2(n22539), .B1(n22957), .B2(n22538), .O(
        n22655) );
  AOI22S U28094 ( .A1(n22625), .A2(gray_img[353]), .B1(gray_img[865]), .B2(
        n22513), .O(n22545) );
  AOI22S U28095 ( .A1(n22935), .A2(gray_img[1145]), .B1(gray_img[1889]), .B2(
        n22794), .O(n22544) );
  ND2S U28096 ( .I1(n15918), .I2(gray_img[241]), .O(n22543) );
  MOAI1S U28097 ( .A1(n22540), .A2(n25996), .B1(gray_img[1257]), .B2(n22936), 
        .O(n22541) );
  AO12S U28098 ( .B1(gray_img[1657]), .B2(n22694), .A1(n22541), .O(n22542) );
  AN4B1S U28099 ( .I1(n22545), .I2(n22544), .I3(n22543), .B1(n22542), .O(
        n22594) );
  AOI22S U28100 ( .A1(gray_img[1529]), .A2(n21096), .B1(n22837), .B2(
        gray_img[361]), .O(n22550) );
  AOI22S U28101 ( .A1(n22762), .A2(gray_img[489]), .B1(n22847), .B2(
        gray_img[1513]), .O(n22549) );
  ND2S U28102 ( .I1(n22663), .I2(gray_img[1137]), .O(n22548) );
  INV1S U28103 ( .I(gray_img[1393]), .O(n27905) );
  MOAI1S U28104 ( .A1(n22797), .A2(n27905), .B1(n22828), .B2(gray_img[1009]), 
        .O(n22546) );
  AO12S U28105 ( .B1(gray_img[1401]), .B2(n21120), .A1(n22546), .O(n22547) );
  AN4B1S U28106 ( .I1(n22550), .I2(n22549), .I3(n22548), .B1(n22547), .O(
        n22593) );
  MOAI1S U28107 ( .A1(n22882), .A2(intadd_32_CI), .B1(n22657), .B2(
        gray_img[745]), .O(n22552) );
  INV1S U28108 ( .I(gray_img[761]), .O(n26332) );
  MOAI1S U28109 ( .A1(n22803), .A2(n26332), .B1(n22785), .B2(gray_img[377]), 
        .O(n22551) );
  NR2 U28110 ( .I1(n22552), .I2(n22551), .O(n22555) );
  AOI22S U28111 ( .A1(n22802), .A2(gray_img[1001]), .B1(gray_img[617]), .B2(
        n22795), .O(n22554) );
  ND2S U28112 ( .I1(n22863), .I2(gray_img[1905]), .O(n22553) );
  ND3S U28113 ( .I1(n22555), .I2(n22554), .I3(n22553), .O(n22572) );
  ND2S U28114 ( .I1(n22893), .I2(gray_img[97]), .O(n22558) );
  AOI22S U28115 ( .A1(n22619), .A2(gray_img[497]), .B1(gray_img[753]), .B2(
        n22695), .O(n22557) );
  AOI22S U28116 ( .A1(n15921), .A2(gray_img[1265]), .B1(gray_img[1649]), .B2(
        n15919), .O(n22556) );
  ND3S U28117 ( .I1(n22558), .I2(n22557), .I3(n22556), .O(n22571) );
  ND2S U28118 ( .I1(n22664), .I2(gray_img[1521]), .O(n22565) );
  ND2S U28119 ( .I1(n22819), .I2(gray_img[1017]), .O(n22564) );
  ND2S U28120 ( .I1(n22900), .I2(gray_img[105]), .O(n22563) );
  ND2S U28121 ( .I1(n22812), .I2(gray_img[2017]), .O(n22561) );
  AOI22S U28122 ( .A1(gray_img[2033]), .A2(n22679), .B1(gray_img[249]), .B2(
        n21089), .O(n22560) );
  ND2S U28123 ( .I1(gray_img[113]), .I2(n22901), .O(n22559) );
  ND3S U28124 ( .I1(n22561), .I2(n22560), .I3(n22559), .O(n22562) );
  AN4B1S U28125 ( .I1(n22565), .I2(n22564), .I3(n22563), .B1(n22562), .O(
        n22569) );
  AOI22S U28126 ( .A1(n22566), .A2(gray_img[993]), .B1(gray_img[737]), .B2(
        n22909), .O(n22568) );
  AOI22S U28127 ( .A1(n22630), .A2(gray_img[609]), .B1(gray_img[481]), .B2(
        n22686), .O(n22567) );
  ND3S U28128 ( .I1(n22569), .I2(n22568), .I3(n22567), .O(n22570) );
  NR3 U28129 ( .I1(n22572), .I2(n22571), .I3(n22570), .O(n22579) );
  AOI22S U28130 ( .A1(n21090), .A2(gray_img[1273]), .B1(n21137), .B2(
        gray_img[121]), .O(n22578) );
  ND2S U28131 ( .I1(n22755), .I2(gray_img[2041]), .O(n22577) );
  AOI22S U28132 ( .A1(n21152), .A2(gray_img[633]), .B1(gray_img[889]), .B2(
        n22813), .O(n22575) );
  AOI22S U28133 ( .A1(n21155), .A2(gray_img[1129]), .B1(gray_img[1769]), .B2(
        n22921), .O(n22574) );
  AOI22S U28134 ( .A1(n22861), .A2(gray_img[1385]), .B1(gray_img[1897]), .B2(
        n22937), .O(n22573) );
  ND3S U28135 ( .I1(n22575), .I2(n22574), .I3(n22573), .O(n22576) );
  AN4B1S U28136 ( .I1(n22579), .I2(n22578), .I3(n22577), .B1(n22576), .O(
        n22591) );
  AOI22S U28137 ( .A1(n15915), .A2(gray_img[625]), .B1(gray_img[881]), .B2(
        n22930), .O(n22590) );
  AOI22S U28138 ( .A1(n22703), .A2(gray_img[1121]), .B1(gray_img[1641]), .B2(
        n22656), .O(n22583) );
  AOI22S U28139 ( .A1(n22864), .A2(gray_img[1913]), .B1(gray_img[1377]), .B2(
        n22934), .O(n22582) );
  AOI22S U28140 ( .A1(n22836), .A2(gray_img[233]), .B1(gray_img[873]), .B2(
        n22932), .O(n22581) );
  MOAI1S U28141 ( .A1(n22670), .A2(intadd_36_CI), .B1(n22610), .B2(
        gray_img[225]), .O(n22580) );
  AN4B1S U28142 ( .I1(n22583), .I2(n22582), .I3(n22581), .B1(n22580), .O(
        n22584) );
  OA12S U28143 ( .B1(intadd_5_CI), .B2(n22853), .A1(n22584), .O(n22589) );
  ND2S U28144 ( .I1(n15905), .I2(gray_img[369]), .O(n22587) );
  AOI22S U28145 ( .A1(n22881), .A2(gray_img[505]), .B1(gray_img[1505]), .B2(
        n21106), .O(n22586) );
  AOI22S U28146 ( .A1(n22770), .A2(gray_img[1761]), .B1(gray_img[1249]), .B2(
        n22838), .O(n22585) );
  ND3S U28147 ( .I1(n22587), .I2(n22586), .I3(n22585), .O(n22588) );
  AN4B1S U28148 ( .I1(n22591), .I2(n22590), .I3(n22589), .B1(n22588), .O(
        n22592) );
  AOI22S U28149 ( .A1(n22727), .A2(gray_img[1865]), .B1(n22894), .B2(
        gray_img[977]), .O(n22599) );
  AOI22S U28150 ( .A1(gray_img[1369]), .A2(n21120), .B1(n22909), .B2(
        gray_img[705]), .O(n22598) );
  ND2S U28151 ( .I1(n22863), .I2(gray_img[1873]), .O(n22597) );
  AOI22S U28152 ( .A1(n22933), .A2(gray_img[201]), .B1(gray_img[1089]), .B2(
        n22703), .O(n22595) );
  OAI12HS U28153 ( .B1(n22797), .B2(intadd_140_CI), .A1(n22595), .O(n22596) );
  AN4B1S U28154 ( .I1(n22599), .I2(n22598), .I3(n22597), .B1(n22596), .O(
        n22651) );
  ND2S U28155 ( .I1(n15915), .I2(gray_img[593]), .O(n22605) );
  AOI22S U28156 ( .A1(n22762), .A2(gray_img[457]), .B1(gray_img[1113]), .B2(
        n22935), .O(n22604) );
  AOI22S U28157 ( .A1(n22837), .A2(gray_img[329]), .B1(gray_img[841]), .B2(
        n22932), .O(n22603) );
  AOI22S U28158 ( .A1(gray_img[849]), .A2(n22930), .B1(n21106), .B2(
        gray_img[1473]), .O(n22600) );
  OAI12HS U28159 ( .B1(n22601), .B2(n25512), .A1(n22600), .O(n22602) );
  AN4B1S U28160 ( .I1(n22605), .I2(n22604), .I3(n22603), .B1(n22602), .O(
        n22650) );
  ND2S U28161 ( .I1(n22931), .I2(gray_img[1993]), .O(n22617) );
  ND2S U28162 ( .I1(n21152), .I2(gray_img[601]), .O(n22609) );
  AOI22S U28163 ( .A1(n22921), .A2(gray_img[1737]), .B1(gray_img[1225]), .B2(
        n22936), .O(n22608) );
  AOI22S U28164 ( .A1(n22934), .A2(gray_img[1345]), .B1(gray_img[1097]), .B2(
        n21155), .O(n22607) );
  MOAI1S U28165 ( .A1(n22875), .A2(intadd_57_CI), .B1(n22656), .B2(
        gray_img[1609]), .O(n22606) );
  AN4B1S U28166 ( .I1(n22609), .I2(n22608), .I3(n22607), .B1(n22606), .O(
        n22616) );
  AOI22S U28167 ( .A1(n15918), .A2(gray_img[209]), .B1(gray_img[337]), .B2(
        n15905), .O(n22615) );
  ND2S U28168 ( .I1(n22663), .I2(gray_img[1105]), .O(n22613) );
  AOI22S U28169 ( .A1(n22513), .A2(gray_img[833]), .B1(gray_img[193]), .B2(
        n22610), .O(n22612) );
  AOI22S U28170 ( .A1(n22864), .A2(gray_img[1881]), .B1(gray_img[1857]), .B2(
        n22794), .O(n22611) );
  ND3S U28171 ( .I1(n22613), .I2(n22612), .I3(n22611), .O(n22614) );
  AN4B1S U28172 ( .I1(n22617), .I2(n22616), .I3(n22615), .B1(n22614), .O(
        n22648) );
  MOAI1S U28173 ( .A1(n22725), .A2(intadd_96_CI), .B1(n21089), .B2(
        gray_img[217]), .O(n22624) );
  INV1S U28174 ( .I(gray_img[1625]), .O(n25525) );
  MOAI1S U28175 ( .A1(n22618), .A2(n25525), .B1(n21096), .B2(gray_img[1497]), 
        .O(n22623) );
  ND2S U28176 ( .I1(n22755), .I2(gray_img[2009]), .O(n22621) );
  AOI22S U28177 ( .A1(n22846), .A2(gray_img[1353]), .B1(n22619), .B2(
        gray_img[465]), .O(n22620) );
  OAI112HS U28178 ( .C1(n22924), .C2(intadd_188_B_0_), .A1(n22621), .B1(n22620), .O(n22622) );
  NR3 U28179 ( .I1(n22624), .I2(n22623), .I3(n22622), .O(n22647) );
  AOI22S U28180 ( .A1(n22735), .A2(gray_img[345]), .B1(gray_img[473]), .B2(
        n22736), .O(n22629) );
  AOI22S U28181 ( .A1(n22770), .A2(gray_img[1729]), .B1(gray_img[321]), .B2(
        n22625), .O(n22628) );
  AOI22S U28182 ( .A1(n22786), .A2(gray_img[1753]), .B1(gray_img[729]), .B2(
        n22883), .O(n22627) );
  MOAI1S U28183 ( .A1(n22670), .A2(intadd_42_CI), .B1(n22838), .B2(
        gray_img[1217]), .O(n22626) );
  AN4B1S U28184 ( .I1(n22629), .I2(n22628), .I3(n22627), .B1(n22626), .O(
        n22641) );
  AOI22S U28185 ( .A1(n22686), .A2(gray_img[449]), .B1(gray_img[969]), .B2(
        n22802), .O(n22640) );
  AOI22S U28186 ( .A1(n22657), .A2(gray_img[713]), .B1(gray_img[585]), .B2(
        n22795), .O(n22639) );
  AOI22S U28187 ( .A1(n22630), .A2(gray_img[577]), .B1(gray_img[961]), .B2(
        n22911), .O(n22637) );
  ND2S U28188 ( .I1(n22900), .I2(gray_img[73]), .O(n22634) );
  ND2S U28189 ( .I1(n22812), .I2(gray_img[1985]), .O(n22633) );
  ND2S U28190 ( .I1(gray_img[81]), .I2(n22901), .O(n22632) );
  INV1S U28191 ( .I(gray_img[1241]), .O(n28289) );
  MOAI1S U28192 ( .A1(n28289), .A2(n22789), .B1(gray_img[2001]), .B2(n22679), 
        .O(n22631) );
  AN4B1S U28193 ( .I1(n22634), .I2(n22633), .I3(n22632), .B1(n22631), .O(
        n22636) );
  ND2S U28194 ( .I1(n22819), .I2(gray_img[985]), .O(n22635) );
  ND3S U28195 ( .I1(n22637), .I2(n22636), .I3(n22635), .O(n22638) );
  AN4B1S U28196 ( .I1(n22641), .I2(n22640), .I3(n22639), .B1(n22638), .O(
        n22646) );
  ND2S U28197 ( .I1(n22893), .I2(gray_img[65]), .O(n22644) );
  AOI22S U28198 ( .A1(n22695), .A2(gray_img[721]), .B1(gray_img[1233]), .B2(
        n15921), .O(n22643) );
  AOI22S U28199 ( .A1(n22796), .A2(gray_img[1745]), .B1(gray_img[1489]), .B2(
        n22664), .O(n22642) );
  ND3S U28200 ( .I1(n22644), .I2(n22643), .I3(n22642), .O(n22645) );
  AN4B1S U28201 ( .I1(n22648), .I2(n22647), .I3(n22646), .B1(n22645), .O(
        n22649) );
  ND3S U28202 ( .I1(n22651), .I2(n22650), .I3(n22649), .O(n22652) );
  AOI22S U28203 ( .A1(n22959), .A2(n22653), .B1(n22782), .B2(n22652), .O(
        n22654) );
  AOI22S U28204 ( .A1(n22934), .A2(gray_img[1285]), .B1(gray_img[1549]), .B2(
        n22656), .O(n22662) );
  AOI22S U28205 ( .A1(n22883), .A2(gray_img[669]), .B1(gray_img[781]), .B2(
        n22932), .O(n22661) );
  AOI22S U28206 ( .A1(n22657), .A2(gray_img[653]), .B1(gray_img[413]), .B2(
        n22881), .O(n22660) );
  MOAI1S U28207 ( .A1(n22658), .A2(n28742), .B1(gray_img[1805]), .B2(n22727), 
        .O(n22659) );
  AN4B1S U28208 ( .I1(n22662), .I2(n22661), .I3(n22660), .B1(n22659), .O(
        n22717) );
  AOI22S U28209 ( .A1(gray_img[541]), .A2(n21152), .B1(n22810), .B2(
        gray_img[645]), .O(n22669) );
  AOI22S U28210 ( .A1(n22837), .A2(gray_img[269]), .B1(n22921), .B2(
        gray_img[1677]), .O(n22668) );
  ND2S U28211 ( .I1(n22663), .I2(gray_img[1045]), .O(n22667) );
  INV1S U28212 ( .I(gray_img[1037]), .O(n26623) );
  MOAI1S U28213 ( .A1(n26623), .A2(n22848), .B1(n22664), .B2(gray_img[1429]), 
        .O(n22665) );
  AO12S U28214 ( .B1(n15918), .B2(gray_img[149]), .A1(n22665), .O(n22666) );
  AN4B1S U28215 ( .I1(n22669), .I2(n22668), .I3(n22667), .B1(n22666), .O(
        n22716) );
  AOI22S U28216 ( .A1(n21106), .A2(gray_img[1413]), .B1(gray_img[1669]), .B2(
        n22770), .O(n22674) );
  AOI22S U28217 ( .A1(n22625), .A2(gray_img[261]), .B1(gray_img[133]), .B2(
        n22610), .O(n22673) );
  AOI22S U28218 ( .A1(n22872), .A2(gray_img[1157]), .B1(gray_img[773]), .B2(
        n22513), .O(n22672) );
  MOAI1S U28219 ( .A1(n22670), .A2(n26596), .B1(n22785), .B2(gray_img[285]), 
        .O(n22671) );
  AN4B1S U28220 ( .I1(n22674), .I2(n22673), .I3(n22672), .B1(n22671), .O(
        n22693) );
  AOI22S U28221 ( .A1(n22795), .A2(gray_img[525]), .B1(gray_img[1693]), .B2(
        n22786), .O(n22678) );
  ND2S U28222 ( .I1(n22863), .I2(gray_img[1813]), .O(n22677) );
  AOI22S U28223 ( .A1(n22911), .A2(gray_img[901]), .B1(gray_img[909]), .B2(
        n22910), .O(n22676) );
  INV1S U28224 ( .I(gray_img[1301]), .O(n29755) );
  NR2 U28225 ( .I1(n29755), .I2(n22797), .O(n22675) );
  AN4B1S U28226 ( .I1(n22678), .I2(n22677), .I3(n22676), .B1(n22675), .O(
        n22692) );
  ND2S U28227 ( .I1(n22893), .I2(gray_img[5]), .O(n22691) );
  AOI22S U28228 ( .A1(n22896), .A2(gray_img[1685]), .B1(gray_img[1557]), .B2(
        n15919), .O(n22689) );
  INV1S U28229 ( .I(gray_img[13]), .O(n23426) );
  NR2 U28230 ( .I1(n23426), .I2(n22811), .O(n22685) );
  INV1S U28231 ( .I(gray_img[157]), .O(n27872) );
  ND2S U28232 ( .I1(n22812), .I2(gray_img[1925]), .O(n22681) );
  AOI22S U28233 ( .A1(gray_img[21]), .A2(n22901), .B1(gray_img[1941]), .B2(
        n22679), .O(n22680) );
  OAI112HS U28234 ( .C1(n21828), .C2(n27872), .A1(n22681), .B1(n22680), .O(
        n22684) );
  INV1S U28235 ( .I(gray_img[925]), .O(n29282) );
  NR2 U28236 ( .I1(n29282), .I2(n22682), .O(n22683) );
  NR3 U28237 ( .I1(n22685), .I2(n22684), .I3(n22683), .O(n22688) );
  AOI22S U28238 ( .A1(n22630), .A2(gray_img[517]), .B1(gray_img[389]), .B2(
        n22686), .O(n22687) );
  ND3S U28239 ( .I1(n22689), .I2(n22688), .I3(n22687), .O(n22690) );
  AN4B1S U28240 ( .I1(n22693), .I2(n22692), .I3(n22691), .B1(n22690), .O(
        n22702) );
  AOI22S U28241 ( .A1(n22694), .A2(gray_img[1565]), .B1(gray_img[1181]), .B2(
        n21090), .O(n22701) );
  ND2S U28242 ( .I1(n22919), .I2(gray_img[1949]), .O(n22700) );
  AOI22S U28243 ( .A1(n21120), .A2(gray_img[1309]), .B1(n21137), .B2(
        gray_img[29]), .O(n22698) );
  AOI22S U28244 ( .A1(n22847), .A2(gray_img[1421]), .B1(n22828), .B2(
        gray_img[917]), .O(n22697) );
  AOI22S U28245 ( .A1(n22695), .A2(gray_img[661]), .B1(gray_img[1173]), .B2(
        n15921), .O(n22696) );
  ND3S U28246 ( .I1(n22698), .I2(n22697), .I3(n22696), .O(n22699) );
  AN4B1S U28247 ( .I1(n22702), .I2(n22701), .I3(n22700), .B1(n22699), .O(
        n22714) );
  AOI22S U28248 ( .A1(n15915), .A2(gray_img[533]), .B1(gray_img[789]), .B2(
        n22930), .O(n22713) );
  AOI22S U28249 ( .A1(n22813), .A2(gray_img[797]), .B1(gray_img[1437]), .B2(
        n21096), .O(n22707) );
  AOI22S U28250 ( .A1(n22794), .A2(gray_img[1797]), .B1(gray_img[1029]), .B2(
        n22703), .O(n22706) );
  AOI22S U28251 ( .A1(n22846), .A2(gray_img[1293]), .B1(gray_img[1165]), .B2(
        n22936), .O(n22705) );
  INV1S U28252 ( .I(gray_img[1933]), .O(n29408) );
  NR2 U28253 ( .I1(n29408), .I2(n22853), .O(n22704) );
  AN4B1S U28254 ( .I1(n22707), .I2(n22706), .I3(n22705), .B1(n22704), .O(
        n22712) );
  ND2S U28255 ( .I1(n15905), .I2(gray_img[277]), .O(n22710) );
  AOI22S U28256 ( .A1(n22933), .A2(gray_img[141]), .B1(gray_img[397]), .B2(
        n22862), .O(n22709) );
  AOI22S U28257 ( .A1(n22935), .A2(gray_img[1053]), .B1(gray_img[1821]), .B2(
        n22787), .O(n22708) );
  ND3S U28258 ( .I1(n22710), .I2(n22709), .I3(n22708), .O(n22711) );
  AN4B1S U28259 ( .I1(n22714), .I2(n22713), .I3(n22712), .B1(n22711), .O(
        n22715) );
  AOI22S U28260 ( .A1(n22895), .A2(gray_img[469]), .B1(gray_img[1621]), .B2(
        n15919), .O(n22723) );
  AOI22S U28261 ( .A1(n22936), .A2(gray_img[1229]), .B1(n22920), .B2(
        gray_img[725]), .O(n22722) );
  ND2S U28262 ( .I1(n21096), .I2(gray_img[1501]), .O(n22721) );
  INV1S U28263 ( .I(gray_img[1477]), .O(n23508) );
  MOAI1S U28264 ( .A1(n22718), .A2(n23508), .B1(gray_img[1373]), .B2(n21120), 
        .O(n22719) );
  AO12S U28265 ( .B1(gray_img[1877]), .B2(n22863), .A1(n22719), .O(n22720) );
  AN4B1S U28266 ( .I1(n22723), .I2(n22722), .I3(n22721), .B1(n22720), .O(
        n22780) );
  ND2S U28267 ( .I1(n22929), .I2(gray_img[1109]), .O(n22731) );
  AOI22S U28268 ( .A1(n22724), .A2(gray_img[845]), .B1(n21155), .B2(
        gray_img[1101]), .O(n22730) );
  AOI22S U28269 ( .A1(n22810), .A2(gray_img[709]), .B1(gray_img[973]), .B2(
        n22910), .O(n22729) );
  INV1S U28270 ( .I(gray_img[861]), .O(n23074) );
  MOAI1S U28271 ( .A1(n22725), .A2(n23074), .B1(n22686), .B2(gray_img[453]), 
        .O(n22726) );
  AO12S U28272 ( .B1(gray_img[1869]), .B2(n22727), .A1(n22726), .O(n22728) );
  AN4B1S U28273 ( .I1(n22731), .I2(n22730), .I3(n22729), .B1(n22728), .O(
        n22779) );
  ND2S U28274 ( .I1(n22893), .I2(gray_img[69]), .O(n22734) );
  AOI22S U28275 ( .A1(n22828), .A2(gray_img[981]), .B1(gray_img[1749]), .B2(
        n22896), .O(n22733) );
  ND2S U28276 ( .I1(n21137), .I2(gray_img[93]), .O(n22732) );
  ND3S U28277 ( .I1(n22734), .I2(n22733), .I3(n22732), .O(n22761) );
  AOI22S U28278 ( .A1(n22786), .A2(gray_img[1757]), .B1(gray_img[349]), .B2(
        n22735), .O(n22740) );
  AOI22S U28279 ( .A1(n22883), .A2(gray_img[733]), .B1(gray_img[477]), .B2(
        n22736), .O(n22739) );
  AOI22S U28280 ( .A1(n22888), .A2(gray_img[717]), .B1(gray_img[589]), .B2(
        n22795), .O(n22738) );
  INV1S U28281 ( .I(gray_img[1365]), .O(n28380) );
  NR2 U28282 ( .I1(n28380), .I2(n22797), .O(n22737) );
  AN4B1S U28283 ( .I1(n22740), .I2(n22739), .I3(n22738), .B1(n22737), .O(
        n22749) );
  AOI22S U28284 ( .A1(n22630), .A2(gray_img[581]), .B1(gray_img[965]), .B2(
        n22911), .O(n22746) );
  ND2S U28285 ( .I1(n22819), .I2(gray_img[989]), .O(n22745) );
  ND2S U28286 ( .I1(n22812), .I2(gray_img[1989]), .O(n22744) );
  INV1S U28287 ( .I(gray_img[77]), .O(n23597) );
  AOI22S U28288 ( .A1(gray_img[2005]), .A2(n22679), .B1(gray_img[597]), .B2(
        n15915), .O(n22742) );
  AOI22S U28289 ( .A1(gray_img[1245]), .A2(n21090), .B1(gray_img[85]), .B2(
        n22901), .O(n22741) );
  OAI112HS U28290 ( .C1(n22811), .C2(n23597), .A1(n22742), .B1(n22741), .O(
        n22743) );
  AN4B1S U28291 ( .I1(n22746), .I2(n22745), .I3(n22744), .B1(n22743), .O(
        n22748) );
  AOI22S U28292 ( .A1(n22664), .A2(gray_img[1493]), .B1(gray_img[1237]), .B2(
        n15921), .O(n22747) );
  ND3S U28293 ( .I1(n22749), .I2(n22748), .I3(n22747), .O(n22760) );
  AOI22S U28294 ( .A1(n22874), .A2(gray_img[1613]), .B1(gray_img[1741]), .B2(
        n22921), .O(n22754) );
  AOI22S U28295 ( .A1(n22846), .A2(gray_img[1357]), .B1(gray_img[1485]), .B2(
        n22847), .O(n22753) );
  AOI22S U28296 ( .A1(n22934), .A2(gray_img[1349]), .B1(gray_img[1093]), .B2(
        n22703), .O(n22752) );
  INV1S U28297 ( .I(gray_img[605]), .O(n27033) );
  NR2 U28298 ( .I1(n27033), .I2(n22750), .O(n22751) );
  AN4B1S U28299 ( .I1(n22754), .I2(n22753), .I3(n22752), .B1(n22751), .O(
        n22758) );
  AOI22S U28300 ( .A1(n21089), .A2(gray_img[221]), .B1(gray_img[1629]), .B2(
        n22918), .O(n22757) );
  ND2S U28301 ( .I1(n22755), .I2(gray_img[2013]), .O(n22756) );
  ND3S U28302 ( .I1(n22758), .I2(n22757), .I3(n22756), .O(n22759) );
  NR3 U28303 ( .I1(n22761), .I2(n22760), .I3(n22759), .O(n22777) );
  ND2S U28304 ( .I1(n22931), .I2(gray_img[1997]), .O(n22768) );
  AOI22S U28305 ( .A1(n22625), .A2(gray_img[325]), .B1(gray_img[837]), .B2(
        n22513), .O(n22767) );
  AOI22S U28306 ( .A1(n22837), .A2(gray_img[333]), .B1(gray_img[205]), .B2(
        n22933), .O(n22766) );
  AOI22S U28307 ( .A1(n22935), .A2(gray_img[1117]), .B1(gray_img[1861]), .B2(
        n22794), .O(n22764) );
  AOI22S U28308 ( .A1(n22762), .A2(gray_img[461]), .B1(gray_img[1885]), .B2(
        n22787), .O(n22763) );
  ND2S U28309 ( .I1(n22764), .I2(n22763), .O(n22765) );
  AN4B1S U28310 ( .I1(n22768), .I2(n22767), .I3(n22766), .B1(n22765), .O(
        n22776) );
  AOI22S U28311 ( .A1(n15905), .A2(gray_img[341]), .B1(gray_img[853]), .B2(
        n22930), .O(n22775) );
  ND2S U28312 ( .I1(n15918), .I2(gray_img[213]), .O(n22773) );
  AOI22S U28313 ( .A1(n22770), .A2(gray_img[1733]), .B1(gray_img[1605]), .B2(
        n21097), .O(n22772) );
  AOI22S U28314 ( .A1(n22872), .A2(gray_img[1221]), .B1(gray_img[197]), .B2(
        n22610), .O(n22771) );
  ND3S U28315 ( .I1(n22773), .I2(n22772), .I3(n22771), .O(n22774) );
  AN4B1S U28316 ( .I1(n22777), .I2(n22776), .I3(n22775), .B1(n22774), .O(
        n22778) );
  ND3S U28317 ( .I1(n22780), .I2(n22779), .I3(n22778), .O(n22781) );
  AOI22S U28318 ( .A1(n22784), .A2(n22783), .B1(n22782), .B2(n22781), .O(
        n22961) );
  ND2S U28319 ( .I1(n15905), .I2(gray_img[373]), .O(n22793) );
  AOI22S U28320 ( .A1(n22786), .A2(gray_img[1789]), .B1(gray_img[381]), .B2(
        n22785), .O(n22792) );
  AOI22S U28321 ( .A1(n22770), .A2(gray_img[1765]), .B1(gray_img[869]), .B2(
        n22513), .O(n22791) );
  INV1S U28322 ( .I(gray_img[1277]), .O(n23319) );
  AOI22S U28323 ( .A1(n22625), .A2(gray_img[357]), .B1(gray_img[1917]), .B2(
        n22787), .O(n22788) );
  OAI12HS U28324 ( .B1(n22789), .B2(n23319), .A1(n22788), .O(n22790) );
  AN4B1S U28325 ( .I1(n22793), .I2(n22792), .I3(n22791), .B1(n22790), .O(
        n22860) );
  AOI22S U28326 ( .A1(n22703), .A2(gray_img[1125]), .B1(n22895), .B2(
        gray_img[501]), .O(n22801) );
  AOI22S U28327 ( .A1(n22932), .A2(gray_img[877]), .B1(gray_img[1893]), .B2(
        n22794), .O(n22800) );
  AOI22S U28328 ( .A1(n22795), .A2(gray_img[621]), .B1(gray_img[229]), .B2(
        n22610), .O(n22799) );
  INV1S U28329 ( .I(gray_img[1397]), .O(n27913) );
  MOAI1S U28330 ( .A1(n22797), .A2(n27913), .B1(n22796), .B2(gray_img[1781]), 
        .O(n22798) );
  AN4B1S U28331 ( .I1(n22801), .I2(n22800), .I3(n22799), .B1(n22798), .O(
        n22859) );
  AOI22S U28332 ( .A1(n15918), .A2(gray_img[245]), .B1(gray_img[629]), .B2(
        n15915), .O(n22808) );
  AOI22S U28333 ( .A1(n22630), .A2(gray_img[613]), .B1(gray_img[485]), .B2(
        n22686), .O(n22807) );
  AOI22S U28334 ( .A1(n22802), .A2(gray_img[1005]), .B1(gray_img[749]), .B2(
        n22888), .O(n22806) );
  MOAI1S U28335 ( .A1(n22803), .A2(n26340), .B1(n22881), .B2(gray_img[509]), 
        .O(n22804) );
  AO12S U28336 ( .B1(gray_img[1909]), .B2(n22863), .A1(n22804), .O(n22805) );
  AN4B1S U28337 ( .I1(n22808), .I2(n22807), .I3(n22806), .B1(n22805), .O(
        n22826) );
  AOI22S U28338 ( .A1(n22664), .A2(gray_img[1525]), .B1(gray_img[1269]), .B2(
        n15921), .O(n22825) );
  ND2S U28339 ( .I1(n22893), .I2(gray_img[101]), .O(n22824) );
  AOI22S U28340 ( .A1(n22911), .A2(gray_img[997]), .B1(gray_img[741]), .B2(
        n22810), .O(n22822) );
  NR2 U28341 ( .I1(n27402), .I2(n22811), .O(n22818) );
  ND2S U28342 ( .I1(n22812), .I2(gray_img[2021]), .O(n22816) );
  AOI22S U28343 ( .A1(gray_img[2037]), .A2(n22679), .B1(gray_img[893]), .B2(
        n22813), .O(n22815) );
  AOI22S U28344 ( .A1(gray_img[117]), .A2(n22901), .B1(gray_img[1405]), .B2(
        n21120), .O(n22814) );
  NR2 U28345 ( .I1(n22818), .I2(n22817), .O(n22821) );
  ND2S U28346 ( .I1(n22819), .I2(gray_img[1021]), .O(n22820) );
  ND3S U28347 ( .I1(n22822), .I2(n22821), .I3(n22820), .O(n22823) );
  AN4B1S U28348 ( .I1(n22826), .I2(n22825), .I3(n22824), .B1(n22823), .O(
        n22835) );
  AOI22S U28349 ( .A1(n21089), .A2(gray_img[253]), .B1(gray_img[1533]), .B2(
        n21096), .O(n22834) );
  ND2S U28350 ( .I1(n22919), .I2(gray_img[2045]), .O(n22833) );
  AOI22S U28351 ( .A1(n22918), .A2(gray_img[1661]), .B1(n21137), .B2(
        gray_img[125]), .O(n22831) );
  AOI22S U28352 ( .A1(n22937), .A2(gray_img[1901]), .B1(n22920), .B2(
        gray_img[757]), .O(n22830) );
  AOI22S U28353 ( .A1(n22828), .A2(gray_img[1013]), .B1(gray_img[1653]), .B2(
        n15919), .O(n22829) );
  ND3S U28354 ( .I1(n22831), .I2(n22830), .I3(n22829), .O(n22832) );
  AN4B1S U28355 ( .I1(n22835), .I2(n22834), .I3(n22833), .B1(n22832), .O(
        n22857) );
  AOI22S U28356 ( .A1(n22837), .A2(gray_img[365]), .B1(gray_img[237]), .B2(
        n22836), .O(n22845) );
  AOI22S U28357 ( .A1(n22935), .A2(gray_img[1149]), .B1(gray_img[1381]), .B2(
        n22934), .O(n22844) );
  ND2S U28358 ( .I1(n22929), .I2(gray_img[1141]), .O(n22843) );
  INV1S U28359 ( .I(gray_img[885]), .O(n26383) );
  AOI22S U28360 ( .A1(n21097), .A2(gray_img[1637]), .B1(gray_img[1253]), .B2(
        n22838), .O(n22840) );
  AOI22S U28361 ( .A1(n21106), .A2(gray_img[1509]), .B1(gray_img[493]), .B2(
        n22862), .O(n22839) );
  OAI112HS U28362 ( .C1(n22841), .C2(n26383), .A1(n22840), .B1(n22839), .O(
        n22842) );
  AN4B1S U28363 ( .I1(n22845), .I2(n22844), .I3(n22843), .B1(n22842), .O(
        n22856) );
  AOI22S U28364 ( .A1(n22921), .A2(gray_img[1773]), .B1(gray_img[1261]), .B2(
        n22936), .O(n22852) );
  ND2S U28365 ( .I1(n21152), .I2(gray_img[637]), .O(n22851) );
  AOI22S U28366 ( .A1(n22874), .A2(gray_img[1645]), .B1(gray_img[1389]), .B2(
        n22846), .O(n22850) );
  INV1S U28367 ( .I(gray_img[1133]), .O(n28051) );
  MOAI1S U28368 ( .A1(n22848), .A2(n28051), .B1(n22847), .B2(gray_img[1517]), 
        .O(n22849) );
  AN4B1S U28369 ( .I1(n22852), .I2(n22851), .I3(n22850), .B1(n22849), .O(
        n22855) );
  INV1S U28370 ( .I(gray_img[2029]), .O(n25856) );
  NR2 U28371 ( .I1(n25856), .I2(n22853), .O(n22854) );
  AN4B1S U28372 ( .I1(n22857), .I2(n22856), .I3(n22855), .B1(n22854), .O(
        n22858) );
  AOI22S U28373 ( .A1(n22861), .A2(gray_img[1325]), .B1(n22827), .B2(
        gray_img[1589]), .O(n22871) );
  AOI22S U28374 ( .A1(n22610), .A2(gray_img[165]), .B1(gray_img[429]), .B2(
        n22862), .O(n22870) );
  ND2S U28375 ( .I1(n22863), .I2(gray_img[1845]), .O(n22869) );
  INV1S U28376 ( .I(gray_img[301]), .O(n27283) );
  MOAI1S U28377 ( .A1(n22865), .A2(n27283), .B1(n22864), .B2(gray_img[1853]), 
        .O(n22866) );
  AO12S U28378 ( .B1(gray_img[829]), .B2(n22867), .A1(n22866), .O(n22868) );
  AN4B1S U28379 ( .I1(n22871), .I2(n22870), .I3(n22869), .B1(n22868), .O(
        n22955) );
  ND2S U28380 ( .I1(n15918), .I2(gray_img[181]), .O(n22880) );
  AOI22S U28381 ( .A1(n22873), .A2(gray_img[957]), .B1(n22872), .B2(
        gray_img[1189]), .O(n22879) );
  AOI22S U28382 ( .A1(n21097), .A2(gray_img[1573]), .B1(n22874), .B2(
        gray_img[1581]), .O(n22878) );
  INV1S U28383 ( .I(gray_img[1453]), .O(n28970) );
  MOAI1S U28384 ( .A1(n22875), .A2(n28970), .B1(n21155), .B2(gray_img[1069]), 
        .O(n22876) );
  AO12S U28385 ( .B1(gray_img[189]), .B2(n21089), .A1(n22876), .O(n22877) );
  AN4B1S U28386 ( .I1(n22880), .I2(n22879), .I3(n22878), .B1(n22877), .O(
        n22954) );
  INV1S U28387 ( .I(gray_img[1725]), .O(n29205) );
  MOAI1S U28388 ( .A1(n22882), .A2(n29205), .B1(n22881), .B2(gray_img[445]), 
        .O(n22886) );
  INV1S U28389 ( .I(gray_img[317]), .O(n26497) );
  MOAI1S U28390 ( .A1(n22884), .A2(n26497), .B1(n22883), .B2(gray_img[701]), 
        .O(n22885) );
  NR2 U28391 ( .I1(n22886), .I2(n22885), .O(n22892) );
  AOI22S U28392 ( .A1(n22888), .A2(gray_img[685]), .B1(gray_img[557]), .B2(
        n22887), .O(n22891) );
  ND2S U28393 ( .I1(n22889), .I2(gray_img[1333]), .O(n22890) );
  ND3S U28394 ( .I1(n22892), .I2(n22891), .I3(n22890), .O(n22917) );
  ND2S U28395 ( .I1(n22893), .I2(gray_img[37]), .O(n22899) );
  AOI22S U28396 ( .A1(n22895), .A2(gray_img[437]), .B1(gray_img[949]), .B2(
        n22894), .O(n22898) );
  AOI22S U28397 ( .A1(n22896), .A2(gray_img[1717]), .B1(gray_img[1461]), .B2(
        n22664), .O(n22897) );
  ND2S U28398 ( .I1(n15921), .I2(gray_img[1205]), .O(n22908) );
  ND2S U28399 ( .I1(n22686), .I2(gray_img[421]), .O(n22907) );
  ND2S U28400 ( .I1(n22900), .I2(gray_img[45]), .O(n22906) );
  INV1S U28401 ( .I(gray_img[1957]), .O(n26664) );
  AOI22S U28402 ( .A1(gray_img[1469]), .A2(n21096), .B1(gray_img[1973]), .B2(
        n22679), .O(n22903) );
  AOI22S U28403 ( .A1(gray_img[53]), .A2(n22901), .B1(gray_img[309]), .B2(
        n15905), .O(n22902) );
  OAI112HS U28404 ( .C1(n22904), .C2(n26664), .A1(n22903), .B1(n22902), .O(
        n22905) );
  AN4B1S U28405 ( .I1(n22908), .I2(n22907), .I3(n22906), .B1(n22905), .O(
        n22914) );
  AOI22S U28406 ( .A1(n22630), .A2(gray_img[549]), .B1(gray_img[677]), .B2(
        n22909), .O(n22913) );
  AOI22S U28407 ( .A1(n22911), .A2(gray_img[933]), .B1(gray_img[941]), .B2(
        n22910), .O(n22912) );
  ND3S U28408 ( .I1(n22914), .I2(n22913), .I3(n22912), .O(n22915) );
  NR3 U28409 ( .I1(n22917), .I2(n22916), .I3(n22915), .O(n22928) );
  AOI22S U28410 ( .A1(n21152), .A2(gray_img[573]), .B1(gray_img[1597]), .B2(
        n22918), .O(n22927) );
  AOI22S U28411 ( .A1(n21090), .A2(gray_img[1213]), .B1(gray_img[1341]), .B2(
        n21120), .O(n22926) );
  INV1S U28412 ( .I(gray_img[61]), .O(n27717) );
  ND2S U28413 ( .I1(n22919), .I2(gray_img[1981]), .O(n22923) );
  AOI22S U28414 ( .A1(n22921), .A2(gray_img[1709]), .B1(n22920), .B2(
        gray_img[693]), .O(n22922) );
  OAI112HS U28415 ( .C1(n22924), .C2(n27717), .A1(n22923), .B1(n22922), .O(
        n22925) );
  AN4B1S U28416 ( .I1(n22928), .I2(n22927), .I3(n22926), .B1(n22925), .O(
        n22952) );
  AOI22S U28417 ( .A1(n22930), .A2(gray_img[821]), .B1(gray_img[1077]), .B2(
        n22929), .O(n22951) );
  ND2S U28418 ( .I1(n22931), .I2(gray_img[1965]), .O(n22944) );
  AOI22S U28419 ( .A1(n22933), .A2(gray_img[173]), .B1(gray_img[813]), .B2(
        n22932), .O(n22943) );
  AOI22S U28420 ( .A1(n22935), .A2(gray_img[1085]), .B1(gray_img[1317]), .B2(
        n22934), .O(n22942) );
  AOI22S U28421 ( .A1(n22937), .A2(gray_img[1837]), .B1(gray_img[1197]), .B2(
        n22936), .O(n22940) );
  AOI22S U28422 ( .A1(n22938), .A2(gray_img[1829]), .B1(gray_img[1061]), .B2(
        n22703), .O(n22939) );
  ND2S U28423 ( .I1(n22940), .I2(n22939), .O(n22941) );
  AN4B1S U28424 ( .I1(n22944), .I2(n22943), .I3(n22942), .B1(n22941), .O(
        n22950) );
  ND2S U28425 ( .I1(n15915), .I2(gray_img[565]), .O(n22948) );
  AOI22S U28426 ( .A1(n21106), .A2(gray_img[1445]), .B1(gray_img[1701]), .B2(
        n22770), .O(n22947) );
  AOI22S U28427 ( .A1(n22625), .A2(gray_img[293]), .B1(gray_img[805]), .B2(
        n22513), .O(n22946) );
  ND3S U28428 ( .I1(n22948), .I2(n22947), .I3(n22946), .O(n22949) );
  AN4B1S U28429 ( .I1(n22952), .I2(n22951), .I3(n22950), .B1(n22949), .O(
        n22953) );
  AOI22S U28430 ( .A1(n22959), .A2(n22958), .B1(n22957), .B2(n22956), .O(
        n22960) );
  INV1S U28431 ( .I(gray_img[966]), .O(n22970) );
  INV1S U28432 ( .I(gray_img[839]), .O(n22969) );
  INV1S U28433 ( .I(gray_img[837]), .O(n22966) );
  FA1S U28434 ( .A(gray_img[961]), .B(gray_img[960]), .CI(intadd_99_CI), .CO(
        n22962) );
  FA1S U28435 ( .A(n22988), .B(gray_img[962]), .CI(n22962), .CO(n22963) );
  FA1S U28436 ( .A(n22986), .B(gray_img[963]), .CI(n22963), .CO(n22964) );
  FA1S U28437 ( .A(n22984), .B(gray_img[964]), .CI(n22964), .CO(n22965) );
  MXL2HS U28438 ( .A(n22971), .B(n22970), .S(n22994), .OB(n22996) );
  INV1S U28439 ( .I(n22996), .O(n27196) );
  FA1S U28440 ( .A(gray_img[841]), .B(gray_img[840]), .CI(intadd_98_CI), .CO(
        n22972) );
  FA1S U28441 ( .A(n22973), .B(gray_img[842]), .CI(n22972), .CO(n22974) );
  FA1S U28442 ( .A(n22975), .B(gray_img[843]), .CI(n22974), .CO(n22976) );
  MXL2HS U28443 ( .A(gray_img[974]), .B(gray_img[846]), .S(n23295), .OB(n22997) );
  INV1S U28444 ( .I(n22997), .O(n27193) );
  INV1S U28445 ( .I(gray_img[964]), .O(n22983) );
  INV1S U28446 ( .I(gray_img[963]), .O(n22985) );
  INV1S U28447 ( .I(gray_img[962]), .O(n22987) );
  INV1S U28448 ( .I(gray_img[961]), .O(n22989) );
  MXL2HS U28449 ( .A(gray_img[837]), .B(gray_img[965]), .S(n22994), .OB(n23008) );
  INV1S U28450 ( .I(gray_img[845]), .O(n27178) );
  MXL2HS U28451 ( .A(n27175), .B(n27178), .S(n23295), .OB(n23005) );
  AOI22S U28452 ( .A1(n27196), .A2(n27193), .B1(n22999), .B2(n22998), .O(
        n23002) );
  INV1S U28453 ( .I(n27222), .O(n27224) );
  OAI112HS U28454 ( .C1(n27230), .C2(n23008), .A1(n23007), .B1(n23006), .O(
        n14120) );
  MAO222S U28455 ( .A1(n23010), .B1(gray_img[1058]), .C1(n23009), .O(n23011)
         );
  MXL2HS U28456 ( .A(gray_img[1186]), .B(gray_img[1058]), .S(n23033), .OB(
        n23048) );
  INV1S U28457 ( .I(gray_img[1198]), .O(n23030) );
  INV1S U28458 ( .I(gray_img[1197]), .O(n23028) );
  INV1S U28459 ( .I(gray_img[1196]), .O(n23026) );
  INV1S U28460 ( .I(gray_img[1195]), .O(n23024) );
  INV1S U28461 ( .I(gray_img[1194]), .O(n23022) );
  MXL2HS U28462 ( .A(gray_img[1190]), .B(gray_img[1062]), .S(n23033), .OB(
        n26144) );
  MXL2HS U28463 ( .A(gray_img[1189]), .B(gray_img[1061]), .S(n23033), .OB(
        n29021) );
  MXL2HS U28464 ( .A(gray_img[1188]), .B(gray_img[1060]), .S(n23033), .OB(
        n29026) );
  MXL2HS U28465 ( .A(gray_img[1187]), .B(gray_img[1059]), .S(n23033), .OB(
        n29031) );
  MXL2HS U28466 ( .A(gray_img[1185]), .B(gray_img[1057]), .S(n23033), .OB(
        n23376) );
  MXL2HS U28467 ( .A(gray_img[1184]), .B(gray_img[1056]), .S(n23033), .OB(
        n29050) );
  OR2 U28468 ( .I1(n29680), .I2(n23042), .O(n29049) );
  INV1S U28469 ( .I(n23042), .O(n23043) );
  INV1S U28470 ( .I(n29044), .O(n29046) );
  OA12S U28471 ( .B1(n29849), .B2(n29046), .A1(n23045), .O(n23046) );
  OAI112HS U28472 ( .C1(n23048), .C2(n29049), .A1(n23047), .B1(n23046), .O(
        n14053) );
  INV1S U28473 ( .I(image[6]), .O(n30338) );
  INV1S U28474 ( .I(image[5]), .O(n30421) );
  INV1S U28475 ( .I(image[4]), .O(n30418) );
  INV1S U28476 ( .I(image[3]), .O(n30417) );
  MAO222 U28477 ( .A1(gray_scale_0[0]), .B1(gray_scale_0[1]), .C1(n30415), .O(
        n23049) );
  MAO222 U28478 ( .A1(n30416), .B1(gray_scale_0[2]), .C1(n23049), .O(n23050)
         );
  FA1 U28479 ( .A(n30418), .B(gray_scale_0[4]), .CI(n23051), .CO(n23052) );
  MOAI1S U28480 ( .A1(n23055), .A2(image[7]), .B1(n30349), .B2(n23054), .O(
        n30422) );
  MOAI1S U28481 ( .A1(n30338), .A2(n30420), .B1(gray_scale_0[6]), .B2(n30419), 
        .O(n15738) );
  INV1S U28482 ( .I(gray_img[854]), .O(n23064) );
  INV1S U28483 ( .I(gray_img[853]), .O(n23062) );
  INV1S U28484 ( .I(gray_img[852]), .O(n23060) );
  INV1S U28485 ( .I(gray_img[851]), .O(n23058) );
  MAO222S U28486 ( .A1(gray_img[977]), .B1(gray_img[976]), .C1(intadd_97_CI), 
        .O(n23056) );
  FA1S U28487 ( .A(intadd_97_B_1_), .B(gray_img[978]), .CI(n23056), .CO(n23057) );
  FA1S U28488 ( .A(n23058), .B(gray_img[979]), .CI(n23057), .CO(n23059) );
  FA1S U28489 ( .A(n23060), .B(gray_img[980]), .CI(n23059), .CO(n23061) );
  MXL2HS U28490 ( .A(gray_img[848]), .B(gray_img[976]), .S(n23079), .OB(n23094) );
  INV1S U28491 ( .I(gray_img[991]), .O(n23067) );
  INV1S U28492 ( .I(gray_img[863]), .O(n23078) );
  ND2S U28493 ( .I1(n23067), .I2(n23078), .O(n25148) );
  NR2 U28494 ( .I1(gray_img[855]), .I2(gray_img[983]), .O(n25149) );
  INV1S U28495 ( .I(gray_img[859]), .O(n23070) );
  FA1S U28496 ( .A(gray_img[985]), .B(gray_img[984]), .CI(intadd_96_CI), .CO(
        n23068) );
  FA1S U28497 ( .A(intadd_96_B_1_), .B(gray_img[986]), .CI(n23068), .CO(n23069) );
  FA1S U28498 ( .A(n23070), .B(gray_img[987]), .CI(n23069), .CO(n23071) );
  MXL2HS U28499 ( .A(gray_img[854]), .B(gray_img[982]), .S(n23079), .OB(n23119) );
  MXL2HS U28500 ( .A(gray_img[853]), .B(gray_img[981]), .S(n23079), .OB(n23114) );
  MXL2HS U28501 ( .A(gray_img[852]), .B(gray_img[980]), .S(n23079), .OB(n23109) );
  MXL2HS U28502 ( .A(gray_img[851]), .B(gray_img[979]), .S(n23079), .OB(n23104) );
  MXL2HS U28503 ( .A(gray_img[850]), .B(gray_img[978]), .S(n23079), .OB(n23099) );
  MXL2HS U28504 ( .A(gray_img[849]), .B(gray_img[977]), .S(n23079), .OB(n23127) );
  MUX2S U28505 ( .A(gray_img[856]), .B(gray_img[984]), .S(n23088), .O(n23089)
         );
  AOI22S U28506 ( .A1(n25372), .A2(n25245), .B1(n25370), .B2(n25244), .O(
        n23090) );
  INV1S U28507 ( .I(n25151), .O(n23123) );
  MUX2S U28508 ( .A(n30005), .B(n25151), .S(gray_img[424]), .O(n23091) );
  OA12S U28509 ( .B1(n29734), .B2(n23123), .A1(n23091), .O(n23092) );
  OAI112HS U28510 ( .C1(n23094), .C2(n23126), .A1(n23093), .B1(n23092), .O(
        n13773) );
  OA12S U28511 ( .B1(n29849), .B2(n23123), .A1(n23096), .O(n23097) );
  OAI112HS U28512 ( .C1(n23099), .C2(n23126), .A1(n23098), .B1(n23097), .O(
        n14114) );
  OA12S U28513 ( .B1(n29843), .B2(n23123), .A1(n23101), .O(n23102) );
  OAI112HS U28514 ( .C1(n23104), .C2(n23126), .A1(n23103), .B1(n23102), .O(
        n14113) );
  OA12S U28515 ( .B1(n29837), .B2(n23123), .A1(n23106), .O(n23107) );
  OAI112HS U28516 ( .C1(n23109), .C2(n23126), .A1(n23108), .B1(n23107), .O(
        n14112) );
  OA12S U28517 ( .B1(n29831), .B2(n23123), .A1(n23111), .O(n23112) );
  OAI112HS U28518 ( .C1(n23114), .C2(n23126), .A1(n23113), .B1(n23112), .O(
        n14111) );
  MUX2S U28519 ( .A(n29032), .B(n25151), .S(gray_img[430]), .O(n23116) );
  OA12S U28520 ( .B1(n29825), .B2(n23123), .A1(n23116), .O(n23117) );
  OAI112HS U28521 ( .C1(n23119), .C2(n23126), .A1(n23118), .B1(n23117), .O(
        n14110) );
  OA12S U28522 ( .B1(n29884), .B2(n23123), .A1(n23122), .O(n23124) );
  OAI112HS U28523 ( .C1(n23127), .C2(n23126), .A1(n23125), .B1(n23124), .O(
        n14115) );
  INV1S U28524 ( .I(gray_img[1982]), .O(n23136) );
  INV1S U28525 ( .I(gray_img[1981]), .O(n23134) );
  INV1S U28526 ( .I(gray_img[1980]), .O(n23132) );
  MAO222S U28527 ( .A1(gray_img[1849]), .B1(gray_img[1848]), .C1(intadd_159_CI), .O(n23128) );
  MXL2HS U28528 ( .A(gray_img[1976]), .B(gray_img[1848]), .S(n23151), .OB(
        n23167) );
  INV1S U28529 ( .I(gray_img[1974]), .O(n23148) );
  INV1S U28530 ( .I(gray_img[1973]), .O(n23146) );
  INV1S U28531 ( .I(gray_img[1972]), .O(n23144) );
  INV1S U28532 ( .I(gray_img[1971]), .O(n23142) );
  INV1S U28533 ( .I(gray_img[1970]), .O(n23140) );
  MXL2HS U28534 ( .A(gray_img[1982]), .B(gray_img[1854]), .S(n23151), .OB(
        n23192) );
  MXL2HS U28535 ( .A(gray_img[1981]), .B(gray_img[1853]), .S(n23151), .OB(
        n23187) );
  MXL2HS U28536 ( .A(gray_img[1980]), .B(gray_img[1852]), .S(n23151), .OB(
        n23182) );
  MXL2HS U28537 ( .A(gray_img[1979]), .B(gray_img[1851]), .S(n23151), .OB(
        n23172) );
  MUX2S U28538 ( .A(gray_img[1970]), .B(gray_img[1842]), .S(n23162), .O(n23173) );
  MXL2HS U28539 ( .A(gray_img[1978]), .B(gray_img[1850]), .S(n23151), .OB(
        n23177) );
  MXL2HS U28540 ( .A(gray_img[1977]), .B(gray_img[1849]), .S(n23151), .OB(
        n23201) );
  MUX2S U28541 ( .A(gray_img[1969]), .B(gray_img[1841]), .S(n23162), .O(n23193) );
  OR2 U28542 ( .I1(n29680), .I2(n23160), .O(n23200) );
  INV1S U28543 ( .I(n23160), .O(n23161) );
  MUX2S U28544 ( .A(gray_img[1968]), .B(gray_img[1840]), .S(n23162), .O(n23163) );
  ND2S U28545 ( .I1(n23194), .I2(n23163), .O(n23166) );
  INV1S U28546 ( .I(n23195), .O(n23197) );
  MUX2S U28547 ( .A(n29032), .B(n23195), .S(gray_img[920]), .O(n23164) );
  OA12S U28548 ( .B1(n29734), .B2(n23197), .A1(n23164), .O(n23165) );
  OAI112HS U28549 ( .C1(n23167), .C2(n23200), .A1(n23166), .B1(n23165), .O(
        n13711) );
  ND2S U28550 ( .I1(n23194), .I2(n23168), .O(n23171) );
  OA12S U28551 ( .B1(n29843), .B2(n23197), .A1(n23169), .O(n23170) );
  OAI112HS U28552 ( .C1(n23172), .C2(n23200), .A1(n23171), .B1(n23170), .O(
        n13639) );
  ND2S U28553 ( .I1(n23194), .I2(n23173), .O(n23176) );
  OA12S U28554 ( .B1(n29849), .B2(n23197), .A1(n23174), .O(n23175) );
  OAI112HS U28555 ( .C1(n23177), .C2(n23200), .A1(n23176), .B1(n23175), .O(
        n13660) );
  ND2S U28556 ( .I1(n23194), .I2(n23178), .O(n23181) );
  MUX2S U28557 ( .A(n30005), .B(n23195), .S(gray_img[924]), .O(n23179) );
  OA12S U28558 ( .B1(n29837), .B2(n23197), .A1(n23179), .O(n23180) );
  OAI112HS U28559 ( .C1(n23182), .C2(n23200), .A1(n23181), .B1(n23180), .O(
        n13629) );
  ND2S U28560 ( .I1(n23194), .I2(n23183), .O(n23186) );
  MUX2S U28561 ( .A(n30005), .B(n23195), .S(gray_img[925]), .O(n23184) );
  OA12S U28562 ( .B1(n29831), .B2(n23197), .A1(n23184), .O(n23185) );
  OAI112HS U28563 ( .C1(n23187), .C2(n23200), .A1(n23186), .B1(n23185), .O(
        n15073) );
  ND2S U28564 ( .I1(n23194), .I2(n23188), .O(n23191) );
  MUX2S U28565 ( .A(n30005), .B(n23195), .S(gray_img[926]), .O(n23189) );
  OA12S U28566 ( .B1(n29825), .B2(n23197), .A1(n23189), .O(n23190) );
  OAI112HS U28567 ( .C1(n23192), .C2(n23200), .A1(n23191), .B1(n23190), .O(
        n13825) );
  ND2S U28568 ( .I1(n23194), .I2(n23193), .O(n23199) );
  OA12S U28569 ( .B1(n29884), .B2(n23197), .A1(n23196), .O(n23198) );
  OAI112HS U28570 ( .C1(n23201), .C2(n23200), .A1(n23199), .B1(n23198), .O(
        n13684) );
  INV1S U28571 ( .I(n29350), .O(n23208) );
  INV1S U28572 ( .I(n23202), .O(n23207) );
  OAI12HS U28573 ( .B1(n23208), .B2(n23207), .A1(n23206), .O(n13955) );
  FA1S U28574 ( .A(gray_img[809]), .B(gray_img[808]), .CI(intadd_162_CI), .CO(
        n23209) );
  FA1S U28575 ( .A(n23210), .B(gray_img[810]), .CI(n23209), .CO(n23211) );
  FA1S U28576 ( .A(n23212), .B(gray_img[811]), .CI(n23211), .CO(n23213) );
  MXL2HS U28577 ( .A(gray_img[937]), .B(gray_img[809]), .S(n23232), .OB(n23246) );
  INV1S U28578 ( .I(gray_img[807]), .O(n25023) );
  INV1S U28579 ( .I(gray_img[935]), .O(n25011) );
  ND2S U28580 ( .I1(n25023), .I2(n25011), .O(n25027) );
  NR2 U28581 ( .I1(gray_img[943]), .I2(gray_img[815]), .O(n25028) );
  INV1S U28582 ( .I(gray_img[933]), .O(n23228) );
  INV1S U28583 ( .I(gray_img[932]), .O(n23226) );
  INV1S U28584 ( .I(gray_img[931]), .O(n23224) );
  INV1S U28585 ( .I(gray_img[930]), .O(n23222) );
  MXL2HS U28586 ( .A(gray_img[942]), .B(gray_img[814]), .S(n23232), .OB(n25766) );
  MXL2HS U28587 ( .A(gray_img[941]), .B(gray_img[813]), .S(n23232), .OB(n28689) );
  MXL2HS U28588 ( .A(gray_img[940]), .B(gray_img[812]), .S(n23232), .OB(n28694) );
  MXL2HS U28589 ( .A(gray_img[939]), .B(gray_img[811]), .S(n23232), .OB(n28699) );
  MXL2HS U28590 ( .A(gray_img[938]), .B(gray_img[810]), .S(n23232), .OB(n28704) );
  MXL2HS U28591 ( .A(gray_img[936]), .B(gray_img[808]), .S(n23232), .OB(n28813) );
  OR2 U28592 ( .I1(n29680), .I2(n23239), .O(n28812) );
  AOI22S U28593 ( .A1(n25372), .A2(n25274), .B1(n25370), .B2(n25272), .O(
        n23242) );
  INV1S U28594 ( .I(n28807), .O(n28809) );
  OA12S U28595 ( .B1(n29884), .B2(n28809), .A1(n23243), .O(n23244) );
  OAI112HS U28596 ( .C1(n23246), .C2(n28812), .A1(n23245), .B1(n23244), .O(
        n14270) );
  INV1S U28597 ( .I(gray_img[2015]), .O(n24979) );
  INV1S U28598 ( .I(gray_img[1887]), .O(n24975) );
  ND2S U28599 ( .I1(n24979), .I2(n24975), .O(n24981) );
  NR2 U28600 ( .I1(gray_img[1879]), .I2(gray_img[2007]), .O(n24982) );
  INV1S U28601 ( .I(gray_img[1886]), .O(n23257) );
  INV1S U28602 ( .I(gray_img[1885]), .O(n23255) );
  INV1S U28603 ( .I(gray_img[1884]), .O(n23253) );
  INV1S U28604 ( .I(gray_img[1882]), .O(n23249) );
  FA1S U28605 ( .A(gray_img[2009]), .B(gray_img[2008]), .CI(n23247), .CO(
        n23248) );
  INV1S U28606 ( .I(gray_img[1879]), .O(n23275) );
  INV1S U28607 ( .I(gray_img[2007]), .O(n23273) );
  INV1S U28608 ( .I(gray_img[1877]), .O(n23259) );
  NR2 U28609 ( .I1(gray_img[2005]), .I2(n23259), .O(n23268) );
  INV1S U28610 ( .I(gray_img[2004]), .O(n23266) );
  INV1S U28611 ( .I(gray_img[2003]), .O(n23264) );
  INV1S U28612 ( .I(gray_img[2002]), .O(n23262) );
  INV1S U28613 ( .I(gray_img[2001]), .O(n23260) );
  FA1S U28614 ( .A(gray_img[1873]), .B(gray_img[1872]), .CI(n23260), .CO(
        n23261) );
  FA1S U28615 ( .A(n23262), .B(gray_img[1874]), .CI(n23261), .CO(n23263) );
  NR2 U28616 ( .I1(n23268), .I2(n23267), .O(n23271) );
  INV1S U28617 ( .I(gray_img[2005]), .O(n23269) );
  INV1S U28618 ( .I(gray_img[2006]), .O(n25403) );
  OAI22S U28619 ( .A1(gray_img[1877]), .A2(n23269), .B1(n25403), .B2(
        gray_img[1878]), .O(n23270) );
  MOAI1S U28620 ( .A1(n23271), .A2(n23270), .B1(gray_img[1878]), .B2(n25403), 
        .O(n23272) );
  OAI12HS U28621 ( .B1(gray_img[1879]), .B2(n23273), .A1(n23272), .O(n23274)
         );
  OAI12HS U28622 ( .B1(gray_img[2007]), .B2(n23275), .A1(n23274), .O(n23285)
         );
  MXL2HS U28623 ( .A(gray_img[2006]), .B(gray_img[1878]), .S(n23285), .OB(
        n25480) );
  MXL2HS U28624 ( .A(gray_img[2005]), .B(gray_img[1877]), .S(n23285), .OB(
        n25585) );
  MXL2HS U28625 ( .A(gray_img[2004]), .B(gray_img[1876]), .S(n23285), .OB(
        n25590) );
  MXL2HS U28626 ( .A(gray_img[2003]), .B(gray_img[1875]), .S(n23285), .OB(
        n25595) );
  MXL2HS U28627 ( .A(gray_img[2002]), .B(gray_img[1874]), .S(n23285), .OB(
        n25600) );
  MXL2HS U28628 ( .A(gray_img[2001]), .B(gray_img[1873]), .S(n23285), .OB(
        n25615) );
  INV1S U28629 ( .I(n23284), .O(n23283) );
  NR2 U28630 ( .I1(n29680), .I2(n23283), .O(n25619) );
  OR2 U28631 ( .I1(n29680), .I2(n23284), .O(n25616) );
  INV1S U28632 ( .I(n25616), .O(n23287) );
  MUX2S U28633 ( .A(gray_img[2000]), .B(gray_img[1872]), .S(n23285), .O(n23286) );
  ND2S U28634 ( .I1(n23287), .I2(n23286), .O(n23291) );
  AOI22S U28635 ( .A1(n25217), .A2(n25245), .B1(n25347), .B2(n25244), .O(
        n23288) );
  ND2S U28636 ( .I1(n15888), .I2(n25612), .O(n23289) );
  ND3S U28637 ( .I1(n23291), .I2(n23290), .I3(n23289), .O(n23292) );
  MUX2S U28638 ( .A(gray_img[968]), .B(gray_img[840]), .S(n23295), .O(n23296)
         );
  OAI112HS U28639 ( .C1(n27230), .C2(n23299), .A1(n23298), .B1(n23297), .O(
        n13774) );
  INV1S U28640 ( .I(gray_img[1142]), .O(n23309) );
  INV1S U28641 ( .I(gray_img[1141]), .O(n23307) );
  INV1S U28642 ( .I(gray_img[1140]), .O(n23305) );
  INV1S U28643 ( .I(gray_img[1139]), .O(n23303) );
  INV1S U28644 ( .I(gray_img[1138]), .O(n23301) );
  MXL2HS U28645 ( .A(gray_img[1138]), .B(gray_img[1266]), .S(n23324), .OB(
        n23339) );
  INV1S U28646 ( .I(gray_img[1278]), .O(n23321) );
  INV1S U28647 ( .I(gray_img[1276]), .O(n23317) );
  INV1S U28648 ( .I(gray_img[1275]), .O(n23315) );
  INV1S U28649 ( .I(gray_img[1274]), .O(n23313) );
  FA1S U28650 ( .A(gray_img[1145]), .B(gray_img[1144]), .CI(intadd_68_CI), 
        .CO(n23312) );
  FA1S U28651 ( .A(n23313), .B(gray_img[1146]), .CI(n23312), .CO(n23314) );
  FA1S U28652 ( .A(n23315), .B(gray_img[1147]), .CI(n23314), .CO(n23316) );
  FA1S U28653 ( .A(n23317), .B(gray_img[1148]), .CI(n23316), .CO(n23318) );
  MXL2HS U28654 ( .A(gray_img[1142]), .B(gray_img[1270]), .S(n23324), .OB(
        n23354) );
  MXL2HS U28655 ( .A(gray_img[1141]), .B(gray_img[1269]), .S(n23324), .OB(
        n23344) );
  MXL2HS U28656 ( .A(gray_img[1140]), .B(gray_img[1268]), .S(n23324), .OB(
        n23359) );
  MXL2HS U28657 ( .A(gray_img[1139]), .B(gray_img[1267]), .S(n23324), .OB(
        n23349) );
  MXL2HS U28658 ( .A(gray_img[1137]), .B(gray_img[1265]), .S(n23324), .OB(
        n23371) );
  MXL2HS U28659 ( .A(gray_img[1136]), .B(gray_img[1264]), .S(n23324), .OB(
        n23499) );
  OR2 U28660 ( .I1(n29680), .I2(n23333), .O(n23498) );
  INV1S U28661 ( .I(n23493), .O(n23495) );
  OA12S U28662 ( .B1(n29849), .B2(n23495), .A1(n23336), .O(n23337) );
  OAI112HS U28663 ( .C1(n23339), .C2(n23498), .A1(n23338), .B1(n23337), .O(
        n14008) );
  OA12S U28664 ( .B1(n29831), .B2(n23495), .A1(n23341), .O(n23342) );
  OAI112HS U28665 ( .C1(n23344), .C2(n23498), .A1(n23343), .B1(n23342), .O(
        n14005) );
  OA12S U28666 ( .B1(n29843), .B2(n23495), .A1(n23346), .O(n23347) );
  OAI112HS U28667 ( .C1(n23349), .C2(n23498), .A1(n23348), .B1(n23347), .O(
        n14007) );
  OA12S U28668 ( .B1(n29825), .B2(n23495), .A1(n23351), .O(n23352) );
  OAI112HS U28669 ( .C1(n23354), .C2(n23498), .A1(n23353), .B1(n23352), .O(
        n14004) );
  OA12S U28670 ( .B1(n29837), .B2(n23495), .A1(n23356), .O(n23357) );
  OAI112HS U28671 ( .C1(n23359), .C2(n23498), .A1(n23358), .B1(n23357), .O(
        n14006) );
  MUX2S U28672 ( .A(gray_img[384]), .B(gray_img[256]), .S(n23360), .O(n23361)
         );
  INV1S U28673 ( .I(n30121), .O(n23363) );
  OAI112HS U28674 ( .C1(n23366), .C2(n30125), .A1(n23365), .B1(n23364), .O(
        n13806) );
  OA12S U28675 ( .B1(n29884), .B2(n23495), .A1(n23368), .O(n23369) );
  OAI112HS U28676 ( .C1(n23371), .C2(n23498), .A1(n23370), .B1(n23369), .O(
        n14009) );
  OAI112HS U28677 ( .C1(n23376), .C2(n29049), .A1(n23375), .B1(n23374), .O(
        n14054) );
  INV1S U28678 ( .I(gray_img[455]), .O(n23387) );
  INV1S U28679 ( .I(gray_img[454]), .O(n23385) );
  INV1S U28680 ( .I(gray_img[453]), .O(n23383) );
  INV1S U28681 ( .I(gray_img[452]), .O(n23381) );
  INV1S U28682 ( .I(gray_img[451]), .O(n23379) );
  MAO222S U28683 ( .A1(gray_img[321]), .B1(gray_img[320]), .C1(intadd_120_CI), 
        .O(n23377) );
  FA1S U28684 ( .A(intadd_120_B_1_), .B(gray_img[322]), .CI(n23377), .CO(
        n23378) );
  FA1S U28685 ( .A(n23379), .B(gray_img[323]), .CI(n23378), .CO(n23380) );
  FA1S U28686 ( .A(n23381), .B(gray_img[324]), .CI(n23380), .CO(n23382) );
  FA1S U28687 ( .A(n23383), .B(gray_img[325]), .CI(n23382), .CO(n23384) );
  MXL2HS U28688 ( .A(gray_img[448]), .B(gray_img[320]), .S(n23401), .OB(n23417) );
  INV1S U28689 ( .I(gray_img[335]), .O(n23388) );
  INV1S U28690 ( .I(gray_img[463]), .O(n23400) );
  ND2S U28691 ( .I1(n23388), .I2(n23400), .O(n25249) );
  NR2 U28692 ( .I1(gray_img[455]), .I2(gray_img[327]), .O(n25250) );
  INV1S U28693 ( .I(gray_img[462]), .O(n23398) );
  INV1S U28694 ( .I(gray_img[461]), .O(n23396) );
  INV1S U28695 ( .I(gray_img[460]), .O(n23394) );
  INV1S U28696 ( .I(gray_img[459]), .O(n23392) );
  INV1S U28697 ( .I(gray_img[458]), .O(n23390) );
  FA1S U28698 ( .A(gray_img[329]), .B(gray_img[328]), .CI(intadd_119_CI), .CO(
        n23389) );
  FA1S U28699 ( .A(n23390), .B(gray_img[330]), .CI(n23389), .CO(n23391) );
  MXL2HS U28700 ( .A(gray_img[454]), .B(gray_img[326]), .S(n23401), .OB(n26865) );
  MXL2HS U28701 ( .A(gray_img[453]), .B(gray_img[325]), .S(n23401), .OB(n26906) );
  MXL2HS U28702 ( .A(gray_img[452]), .B(gray_img[324]), .S(n23401), .OB(n26911) );
  MXL2HS U28703 ( .A(gray_img[451]), .B(gray_img[323]), .S(n23401), .OB(n26916) );
  MXL2HS U28704 ( .A(gray_img[450]), .B(gray_img[322]), .S(n23401), .OB(n26921) );
  MXL2HS U28705 ( .A(gray_img[449]), .B(gray_img[321]), .S(n23401), .OB(n26935) );
  OR2 U28706 ( .I1(n29680), .I2(n23408), .O(n26936) );
  INV1S U28707 ( .I(n23408), .O(n23409) );
  MUX2S U28708 ( .A(gray_img[456]), .B(gray_img[328]), .S(n23410), .O(n23411)
         );
  AOI22S U28709 ( .A1(n25246), .A2(n25194), .B1(n25257), .B2(n25193), .O(
        n23412) );
  INV1S U28710 ( .I(n26932), .O(n23414) );
  MUX2S U28711 ( .A(n29032), .B(n26932), .S(gray_img[160]), .O(n23413) );
  OAI112HS U28712 ( .C1(n23417), .C2(n26936), .A1(n23416), .B1(n23415), .O(
        n13804) );
  INV1S U28713 ( .I(gray_img[15]), .O(n23430) );
  FA1S U28714 ( .A(gray_img[137]), .B(gray_img[136]), .CI(n23418), .CO(n23419)
         );
  FA1S U28715 ( .A(n23420), .B(gray_img[138]), .CI(n23419), .CO(n23421) );
  FA1S U28716 ( .A(n23422), .B(gray_img[139]), .CI(n23421), .CO(n23423) );
  FA1S U28717 ( .A(n23424), .B(gray_img[140]), .CI(n23423), .CO(n23425) );
  MXL2HS U28718 ( .A(gray_img[12]), .B(gray_img[140]), .S(n30111), .OB(n23457)
         );
  INV1S U28719 ( .I(gray_img[135]), .O(n23431) );
  INV1S U28720 ( .I(gray_img[7]), .O(n25118) );
  ND2S U28721 ( .I1(n23431), .I2(n25118), .O(n25113) );
  NR2 U28722 ( .I1(gray_img[15]), .I2(gray_img[143]), .O(n25114) );
  INV1S U28723 ( .I(gray_img[6]), .O(n23442) );
  INV1S U28724 ( .I(gray_img[5]), .O(n23440) );
  INV1S U28725 ( .I(gray_img[4]), .O(n23438) );
  INV1S U28726 ( .I(gray_img[2]), .O(n23434) );
  MXL2HS U28727 ( .A(gray_img[14]), .B(gray_img[142]), .S(n30111), .OB(n23477)
         );
  MXL2HS U28728 ( .A(gray_img[13]), .B(gray_img[141]), .S(n30111), .OB(n23472)
         );
  MXL2HS U28729 ( .A(gray_img[11]), .B(gray_img[139]), .S(n30111), .OB(n23462)
         );
  MXL2HS U28730 ( .A(gray_img[10]), .B(gray_img[138]), .S(n30111), .OB(n23467)
         );
  MUX2S U28731 ( .A(gray_img[0]), .B(gray_img[128]), .S(n23444), .O(n30119) );
  MXL2HS U28732 ( .A(gray_img[9]), .B(gray_img[137]), .S(n30111), .OB(n23482)
         );
  OR2 U28733 ( .I1(n29680), .I2(n23450), .O(n30110) );
  AOI22S U28734 ( .A1(n25218), .A2(n25273), .B1(n25216), .B2(n25271), .O(
        n23453) );
  INV1S U28735 ( .I(n30114), .O(n30117) );
  MUX2S U28736 ( .A(n29032), .B(n30114), .S(gray_img[4]), .O(n23454) );
  OA12S U28737 ( .B1(n29837), .B2(n30117), .A1(n23454), .O(n23455) );
  OAI112HS U28738 ( .C1(n23457), .C2(n30110), .A1(n23456), .B1(n23455), .O(
        n14876) );
  MUX2S U28739 ( .A(n30005), .B(n30114), .S(gray_img[3]), .O(n23459) );
  OA12S U28740 ( .B1(n29843), .B2(n30117), .A1(n23459), .O(n23460) );
  OAI112HS U28741 ( .C1(n23462), .C2(n30110), .A1(n23461), .B1(n23460), .O(
        n14677) );
  MUX2S U28742 ( .A(n30005), .B(n30114), .S(gray_img[2]), .O(n23464) );
  OA12S U28743 ( .B1(n29849), .B2(n30117), .A1(n23464), .O(n23465) );
  OAI112HS U28744 ( .C1(n23467), .C2(n30110), .A1(n23466), .B1(n23465), .O(
        n14477) );
  MUX2S U28745 ( .A(n30005), .B(n30114), .S(gray_img[5]), .O(n23469) );
  OA12S U28746 ( .B1(n29831), .B2(n30117), .A1(n23469), .O(n23470) );
  OAI112HS U28747 ( .C1(n23472), .C2(n30110), .A1(n23471), .B1(n23470), .O(
        n15076) );
  MUX2S U28748 ( .A(n29032), .B(n30114), .S(gray_img[6]), .O(n23474) );
  OA12S U28749 ( .B1(n29825), .B2(n30117), .A1(n23474), .O(n23475) );
  OAI112HS U28750 ( .C1(n23477), .C2(n30110), .A1(n23476), .B1(n23475), .O(
        n15465) );
  MUX2S U28751 ( .A(n30005), .B(n30114), .S(gray_img[1]), .O(n23479) );
  OA12S U28752 ( .B1(n29884), .B2(n30117), .A1(n23479), .O(n23480) );
  OAI112HS U28753 ( .C1(n23482), .C2(n30110), .A1(n23481), .B1(n23480), .O(
        n14276) );
  MUX2S U28754 ( .A(gray_img[208]), .B(gray_img[80]), .S(n23483), .O(n23484)
         );
  INV1S U28755 ( .I(n26842), .O(n23486) );
  OAI112HS U28756 ( .C1(n23489), .C2(n26846), .A1(n23488), .B1(n23487), .O(
        n13809) );
  MUX2S U28757 ( .A(gray_img[1272]), .B(gray_img[1144]), .S(n23490), .O(n23491) );
  OA12S U28758 ( .B1(n29734), .B2(n23495), .A1(n23494), .O(n23496) );
  OAI112HS U28759 ( .C1(n23499), .C2(n23498), .A1(n23497), .B1(n23496), .O(
        n13739) );
  INV1S U28760 ( .I(gray_img[1476]), .O(n23506) );
  INV1S U28761 ( .I(gray_img[1475]), .O(n23504) );
  INV1S U28762 ( .I(gray_img[1474]), .O(n23502) );
  INV1S U28763 ( .I(gray_img[1473]), .O(n23500) );
  NR2 U28764 ( .I1(gray_img[1351]), .I2(n23512), .O(n23514) );
  AOI12HS U28765 ( .B1(n23512), .B2(gray_img[1351]), .A1(n23511), .O(n23513)
         );
  MXL2HS U28766 ( .A(gray_img[1472]), .B(gray_img[1344]), .S(n23530), .OB(
        n23543) );
  INV1S U28767 ( .I(gray_img[1359]), .O(n25203) );
  ND2S U28768 ( .I1(n25203), .I2(n25199), .O(n25206) );
  NR2 U28769 ( .I1(gray_img[1351]), .I2(gray_img[1479]), .O(n25207) );
  MXL2HS U28770 ( .A(gray_img[1477]), .B(gray_img[1349]), .S(n23530), .OB(
        n28540) );
  INV1S U28771 ( .I(gray_img[1486]), .O(n23524) );
  INV1S U28772 ( .I(gray_img[1485]), .O(n23522) );
  INV1S U28773 ( .I(gray_img[1484]), .O(n23520) );
  INV1S U28774 ( .I(gray_img[1482]), .O(n23516) );
  MAO222S U28775 ( .A1(gray_img[1353]), .B1(gray_img[1352]), .C1(intadd_57_CI), 
        .O(n23515) );
  MAO222S U28776 ( .A1(n23516), .B1(gray_img[1354]), .C1(n23515), .O(n23517)
         );
  FA1S U28777 ( .A(n23518), .B(gray_img[1355]), .CI(n23517), .CO(n23519) );
  FA1S U28778 ( .A(n23520), .B(gray_img[1356]), .CI(n23519), .CO(n23521) );
  MUX2S U28779 ( .A(gray_img[1484]), .B(gray_img[1356]), .S(n23536), .O(n28547) );
  MXL2HS U28780 ( .A(gray_img[1476]), .B(gray_img[1348]), .S(n23530), .OB(
        n28545) );
  MUX2S U28781 ( .A(gray_img[1483]), .B(gray_img[1355]), .S(n23536), .O(n28552) );
  MXL2HS U28782 ( .A(gray_img[1475]), .B(gray_img[1347]), .S(n23530), .OB(
        n28550) );
  MUX2S U28783 ( .A(gray_img[1482]), .B(gray_img[1354]), .S(n23536), .O(n28557) );
  MXL2HS U28784 ( .A(gray_img[1474]), .B(gray_img[1346]), .S(n23530), .OB(
        n28555) );
  MXL2HS U28785 ( .A(gray_img[1473]), .B(gray_img[1345]), .S(n23530), .OB(
        n28584) );
  MUX2S U28786 ( .A(gray_img[1481]), .B(gray_img[1353]), .S(n23536), .O(n28587) );
  AOI22S U28787 ( .A1(n28540), .A2(n28542), .B1(n23529), .B2(n15976), .O(
        n23532) );
  MXL2HS U28788 ( .A(gray_img[1478]), .B(gray_img[1350]), .S(n23530), .OB(
        n23548) );
  INV1S U28789 ( .I(n23534), .O(n23535) );
  MUX2S U28790 ( .A(gray_img[1480]), .B(gray_img[1352]), .S(n23536), .O(n23537) );
  ND2S U28791 ( .I1(n28588), .I2(n23537), .O(n23542) );
  AOI22S U28792 ( .A1(n25308), .A2(n25194), .B1(n25340), .B2(n25193), .O(
        n23538) );
  INV1S U28793 ( .I(n28581), .O(n23540) );
  OA12S U28794 ( .B1(n29734), .B2(n23540), .A1(n23539), .O(n23541) );
  OAI112HS U28795 ( .C1(n23543), .C2(n28585), .A1(n23542), .B1(n23541), .O(
        n13726) );
  ND2S U28796 ( .I1(n28588), .I2(n23544), .O(n23547) );
  OA12S U28797 ( .B1(gray_img[678]), .B2(n29427), .A1(n28581), .O(n23545) );
  MOAI1S U28798 ( .A1(n28581), .A2(gray_img[678]), .B1(n29825), .B2(n23545), 
        .O(n23546) );
  OAI112HS U28799 ( .C1(n23548), .C2(n28585), .A1(n23547), .B1(n23546), .O(
        n13945) );
  FA1S U28800 ( .A(intadd_25_B_0_), .B(intadd_25_A_0_), .CI(gray_img[1857]), 
        .CO(n23549) );
  FA1S U28801 ( .A(gray_img[1858]), .B(n23550), .CI(n23549), .CO(n23551) );
  FA1S U28802 ( .A(gray_img[1859]), .B(n23552), .CI(n23551), .CO(n23553) );
  MXL2HS U28803 ( .A(gray_img[1984]), .B(gray_img[1856]), .S(n23573), .OB(
        n23589) );
  INV1S U28804 ( .I(gray_img[1871]), .O(n25004) );
  ND2S U28805 ( .I1(n25004), .I2(n25001), .O(n25007) );
  NR2 U28806 ( .I1(gray_img[1991]), .I2(gray_img[1863]), .O(n25008) );
  FA1S U28807 ( .A(gray_img[1865]), .B(gray_img[1864]), .CI(n23561), .CO(
        n23562) );
  FA1S U28808 ( .A(n23563), .B(gray_img[1866]), .CI(n23562), .CO(n23564) );
  FA1S U28809 ( .A(n23565), .B(gray_img[1867]), .CI(n23564), .CO(n23566) );
  MXL2HS U28810 ( .A(gray_img[1990]), .B(gray_img[1862]), .S(n23573), .OB(
        n25635) );
  MXL2HS U28811 ( .A(gray_img[1989]), .B(gray_img[1861]), .S(n23573), .OB(
        n25722) );
  MXL2HS U28812 ( .A(gray_img[1988]), .B(gray_img[1860]), .S(n23573), .OB(
        n25727) );
  MXL2HS U28813 ( .A(gray_img[1987]), .B(gray_img[1859]), .S(n23573), .OB(
        n25732) );
  MXL2HS U28814 ( .A(gray_img[1986]), .B(gray_img[1858]), .S(n23573), .OB(
        n25737) );
  MXL2HS U28815 ( .A(gray_img[1985]), .B(gray_img[1857]), .S(n23573), .OB(
        n25754) );
  MAO222 U28816 ( .A1(n23589), .B1(n25754), .C1(n25757), .O(n23574) );
  MAO222 U28817 ( .A1(n25739), .B1(n25737), .C1(n23574), .O(n23575) );
  FA1S U28818 ( .A(n25734), .B(n25732), .CI(n23575), .CO(n23576) );
  OR2 U28819 ( .I1(n29680), .I2(n23580), .O(n25755) );
  INV1S U28820 ( .I(n23580), .O(n23581) );
  MUX2S U28821 ( .A(gray_img[1992]), .B(gray_img[1864]), .S(n23582), .O(n23583) );
  AOI22S U28822 ( .A1(n25194), .A2(n25217), .B1(n25193), .B2(n25347), .O(
        n23584) );
  INV1S U28823 ( .I(n25751), .O(n23586) );
  OAI112HS U28824 ( .C1(n23589), .C2(n25755), .A1(n23588), .B1(n23587), .O(
        n13710) );
  INV1S U28825 ( .I(gray_img[76]), .O(n23595) );
  FA1S U28826 ( .A(intadd_130_B_0_), .B(intadd_130_A_0_), .CI(gray_img[201]), 
        .CO(n23590) );
  FA1S U28827 ( .A(gray_img[202]), .B(n23591), .CI(n23590), .CO(n23592) );
  FA1S U28828 ( .A(gray_img[203]), .B(n23593), .CI(n23592), .CO(n23594) );
  MXL2HS U28829 ( .A(gray_img[72]), .B(gray_img[200]), .S(n23615), .OB(n23631)
         );
  ND2S U28830 ( .I1(n23602), .I2(n23614), .O(n25261) );
  NR2 U28831 ( .I1(gray_img[79]), .I2(gray_img[207]), .O(n25262) );
  INV1S U28832 ( .I(gray_img[198]), .O(n23612) );
  INV1S U28833 ( .I(gray_img[197]), .O(n23610) );
  INV1S U28834 ( .I(gray_img[196]), .O(n23608) );
  INV1S U28835 ( .I(gray_img[195]), .O(n23606) );
  INV1S U28836 ( .I(gray_img[194]), .O(n23604) );
  FA1S U28837 ( .A(gray_img[65]), .B(gray_img[64]), .CI(intadd_129_CI), .CO(
        n23603) );
  MAO222S U28838 ( .A1(n23604), .B1(gray_img[66]), .C1(n23603), .O(n23605) );
  FA1S U28839 ( .A(n23606), .B(gray_img[67]), .CI(n23605), .CO(n23607) );
  FA1S U28840 ( .A(n23608), .B(gray_img[68]), .CI(n23607), .CO(n23609) );
  MXL2HS U28841 ( .A(gray_img[78]), .B(gray_img[206]), .S(n23615), .OB(n23636)
         );
  MXL2HS U28842 ( .A(gray_img[77]), .B(gray_img[205]), .S(n23615), .OB(n26886)
         );
  MXL2HS U28843 ( .A(gray_img[76]), .B(gray_img[204]), .S(n23615), .OB(n26891)
         );
  MXL2HS U28844 ( .A(gray_img[75]), .B(gray_img[203]), .S(n23615), .OB(n26896)
         );
  MXL2HS U28845 ( .A(gray_img[74]), .B(gray_img[202]), .S(n23615), .OB(n26901)
         );
  MXL2HS U28846 ( .A(gray_img[73]), .B(gray_img[201]), .S(n23615), .OB(n26927)
         );
  OR2 U28847 ( .I1(n29680), .I2(n23622), .O(n26928) );
  INV1S U28848 ( .I(n23622), .O(n23623) );
  MUX2S U28849 ( .A(gray_img[192]), .B(gray_img[64]), .S(n23624), .O(n23625)
         );
  AOI22S U28850 ( .A1(n25194), .A2(n25273), .B1(n25193), .B2(n25271), .O(
        n23626) );
  INV1S U28851 ( .I(n26924), .O(n23628) );
  OAI112HS U28852 ( .C1(n23631), .C2(n26928), .A1(n23630), .B1(n23629), .O(
        n13810) );
  OA12S U28853 ( .B1(gray_img[38]), .B2(n29427), .A1(n26924), .O(n23633) );
  MOAI1S U28854 ( .A1(n26924), .A2(gray_img[38]), .B1(n29825), .B2(n23633), 
        .O(n23634) );
  OAI112HS U28855 ( .C1(n23636), .C2(n26928), .A1(n23635), .B1(n23634), .O(
        n14251) );
  INV1S U28856 ( .I(mem_data_out_reg_shift_1[30]), .O(n23640) );
  AO12T U28857 ( .B1(n24069), .B2(medfilt_state[0]), .A1(medfilt_state[3]), 
        .O(n23984) );
  INV1S U28858 ( .I(n24928), .O(n23639) );
  ND2S U28859 ( .I1(n23637), .I2(medfilt_state[0]), .O(n23638) );
  ND3HT U28860 ( .I1(n24118), .I2(n23639), .I3(n23638), .O(n23782) );
  NR2T U28861 ( .I1(n23984), .I2(n23782), .O(n23687) );
  NR2 U28862 ( .I1(n23640), .I2(n23687), .O(n23674) );
  INV1S U28863 ( .I(n23674), .O(n23677) );
  INV1S U28864 ( .I(mem_data_out_reg_shift_1[26]), .O(n23641) );
  INV1S U28865 ( .I(n23652), .O(n23648) );
  INV1S U28866 ( .I(mem_data_out_reg_shift_1[25]), .O(n23642) );
  INV1S U28867 ( .I(mem_data_out_reg_shift_1[17]), .O(n24265) );
  NR2P U28868 ( .I1(medfilt_state[0]), .I2(n24919), .O(n23986) );
  BUF4CK U28869 ( .I(n23986), .O(n23784) );
  ND2S U28870 ( .I1(n30453), .I2(medfilt_state[0]), .O(n23643) );
  NR2 U28871 ( .I1(medfilt_state[2]), .I2(n23643), .O(n23987) );
  INV2 U28872 ( .I(n23987), .O(n24067) );
  ND2T U28873 ( .I1(n24067), .I2(n24047), .O(n23783) );
  OR2T U28874 ( .I1(n23784), .I2(n23783), .O(n23689) );
  INV4 U28875 ( .I(n23689), .O(n23672) );
  NR2 U28876 ( .I1(n24265), .I2(n23672), .O(n23644) );
  ND2S U28877 ( .I1(n23645), .I2(n24265), .O(n23646) );
  OAI112HS U28878 ( .C1(mem_data_out_reg_shift_1[18]), .C2(n23648), .A1(n23647), .B1(n23646), .O(n23659) );
  INV1S U28879 ( .I(mem_data_out_reg_shift_1[29]), .O(n23649) );
  NR2 U28880 ( .I1(n30456), .I2(n23672), .O(n23650) );
  INV1S U28881 ( .I(mem_data_out_reg_shift_1[18]), .O(n24292) );
  NR2 U28882 ( .I1(n24292), .I2(n23672), .O(n23651) );
  NR2P U28883 ( .I1(n23652), .I2(n23651), .O(n24290) );
  AOI22S U28884 ( .A1(n24316), .A2(mem_data_out_reg_shift_1[21]), .B1(
        mem_data_out_reg_shift_1[18]), .B2(n24290), .O(n23658) );
  INV1S U28885 ( .I(mem_data_out_reg_shift_1[19]), .O(n24283) );
  INV1S U28886 ( .I(mem_data_out_reg_shift_1[27]), .O(n23653) );
  NR2P U28887 ( .I1(n23654), .I2(n15920), .O(n24281) );
  INV1S U28888 ( .I(mem_data_out_reg_shift_1[28]), .O(n23655) );
  NR2T U28889 ( .I1(n23656), .I2(n15906), .O(n24324) );
  AOI22S U28890 ( .A1(n24281), .A2(mem_data_out_reg_shift_1[19]), .B1(
        mem_data_out_reg_shift_1[20]), .B2(n24324), .O(n23657) );
  ND2 U28891 ( .I1(n15920), .I2(n24283), .O(n23664) );
  NR2 U28892 ( .I1(mem_data_out_reg_shift_1[19]), .I2(
        mem_data_out_reg_shift_1[20]), .O(n23660) );
  AOI22S U28893 ( .A1(n15906), .A2(n24327), .B1(n15920), .B2(n23660), .O(
        n23661) );
  OA12S U28894 ( .B1(n24324), .B2(n23664), .A1(n23661), .O(n23671) );
  INV1S U28895 ( .I(n15906), .O(n23663) );
  ND2S U28896 ( .I1(n23664), .I2(n23663), .O(n23669) );
  ND3S U28897 ( .I1(n15920), .I2(n30456), .I3(n24283), .O(n23667) );
  MOAI1 U28898 ( .A1(n24324), .A2(n23667), .B1(n23666), .B2(n30456), .O(n23668) );
  AOI13HS U28899 ( .B1(n30456), .B2(n24327), .B3(n23669), .A1(n23668), .O(
        n23670) );
  OAI12HS U28900 ( .B1(n23671), .B2(n24316), .A1(n23670), .O(n23675) );
  NR2 U28901 ( .I1(n24270), .I2(n23672), .O(n23673) );
  INV2 U28902 ( .I(n23680), .O(n23678) );
  NR2P U28903 ( .I1(mem_data_out_reg_shift_1[23]), .I2(n23678), .O(n23683) );
  INV1S U28904 ( .I(mem_data_out_reg_shift_1[31]), .O(n23679) );
  NR2 U28905 ( .I1(n23679), .I2(n23687), .O(n24601) );
  INV1S U28906 ( .I(n24601), .O(n24342) );
  ND2S U28907 ( .I1(n23689), .I2(mem_data_out_reg_shift_1[23]), .O(n24602) );
  INV1S U28908 ( .I(mem_data_out_reg_shift_1[23]), .O(n24341) );
  NR2F U28909 ( .I1(n23683), .I2(n23682), .O(n23738) );
  ND2P U28910 ( .I1(n23684), .I2(n30242), .O(n24115) );
  NR2T U28911 ( .I1(n24100), .I2(n24115), .O(n23906) );
  INV1S U28912 ( .I(mem_data_out_reg_shift_1[11]), .O(n23802) );
  ND3HT U28913 ( .I1(n24068), .I2(n23993), .I3(n23685), .O(n23863) );
  NR2T U28914 ( .I1(n24069), .I2(n23863), .O(n23905) );
  NR2 U28915 ( .I1(n24285), .I2(n24281), .O(n23694) );
  INV1S U28916 ( .I(mem_data_out_reg_shift_1[10]), .O(n23807) );
  NR2 U28917 ( .I1(n24294), .I2(n24290), .O(n23686) );
  NR2 U28918 ( .I1(n23694), .I2(n23686), .O(n23697) );
  INV1S U28919 ( .I(mem_data_out_reg_shift_1[9]), .O(n23813) );
  OR2T U28920 ( .I1(n23813), .I2(n23905), .O(n23713) );
  OAI12H U28921 ( .B1(n23906), .B2(n24265), .A1(n23713), .O(n24267) );
  INV1S U28922 ( .I(mem_data_out_reg_shift_1[24]), .O(n23688) );
  NR2 U28923 ( .I1(n24267), .I2(n23908), .O(n23691) );
  INV1S U28924 ( .I(n23914), .O(n24566) );
  ND2S U28925 ( .I1(n23908), .I2(n24267), .O(n23690) );
  OAI12HS U28926 ( .B1(n23691), .B2(n24566), .A1(n23690), .O(n23696) );
  ND2S U28927 ( .I1(n24290), .I2(n24294), .O(n23693) );
  ND2S U28928 ( .I1(n24281), .I2(n24285), .O(n23692) );
  OAI12HS U28929 ( .B1(n23694), .B2(n23693), .A1(n23692), .O(n23695) );
  AOI12HS U28930 ( .B1(n23697), .B2(n23696), .A1(n23695), .O(n23712) );
  INV1S U28931 ( .I(mem_data_out_reg_shift_1[13]), .O(n23826) );
  NR2 U28932 ( .I1(n24319), .I2(n24316), .O(n23703) );
  INV1S U28933 ( .I(mem_data_out_reg_shift_1[12]), .O(n23831) );
  OAI12HS U28934 ( .B1(n23906), .B2(n24327), .A1(n23724), .O(n24330) );
  NR2 U28935 ( .I1(n24330), .I2(n24324), .O(n23698) );
  NR2 U28936 ( .I1(n23703), .I2(n23698), .O(n23700) );
  INV1S U28937 ( .I(mem_data_out_reg_shift_1[15]), .O(n23842) );
  OAI12HS U28938 ( .B1(n23906), .B2(n24341), .A1(n24340), .O(n24605) );
  INV1S U28939 ( .I(mem_data_out_reg_shift_1[14]), .O(n23837) );
  OAI12HS U28940 ( .B1(n23906), .B2(n24270), .A1(n23730), .O(n24272) );
  NR2 U28941 ( .I1(n24272), .I2(n24268), .O(n23699) );
  NR2 U28942 ( .I1(n23706), .I2(n23699), .O(n23709) );
  ND2S U28943 ( .I1(n23700), .I2(n23709), .O(n23711) );
  ND2S U28944 ( .I1(n24324), .I2(n24330), .O(n23702) );
  ND2S U28945 ( .I1(n24316), .I2(n24319), .O(n23701) );
  OAI12HS U28946 ( .B1(n23703), .B2(n23702), .A1(n23701), .O(n23708) );
  ND2S U28947 ( .I1(n24268), .I2(n24272), .O(n23705) );
  ND2S U28948 ( .I1(n23956), .I2(n24605), .O(n23704) );
  OAI12HS U28949 ( .B1(n23706), .B2(n23705), .A1(n23704), .O(n23707) );
  AOI12HS U28950 ( .B1(n23709), .B2(n23708), .A1(n23707), .O(n23710) );
  INV1S U28951 ( .I(n24605), .O(n23954) );
  OAI22S U28952 ( .A1(n24283), .A2(n24285), .B1(n24294), .B2(n24292), .O(
        n23721) );
  ND2S U28953 ( .I1(n23714), .I2(n24265), .O(n23715) );
  MOAI1 U28954 ( .A1(n24267), .A2(n24265), .B1(mem_data_out_reg_shift_1[16]), 
        .B2(n23715), .O(n23716) );
  OAI12HS U28955 ( .B1(mem_data_out_reg_shift_1[18]), .B2(n23717), .A1(n23716), 
        .O(n23718) );
  INV1 U28956 ( .I(n23718), .O(n23720) );
  OAI22S U28957 ( .A1(n23721), .A2(n23720), .B1(mem_data_out_reg_shift_1[19]), 
        .B2(n23719), .O(n23722) );
  OAI12HS U28958 ( .B1(n24327), .B2(n24330), .A1(n23722), .O(n23729) );
  INV1S U28959 ( .I(n23723), .O(n23726) );
  INV1S U28960 ( .I(n23724), .O(n23725) );
  AOI22S U28961 ( .A1(n23726), .A2(n30456), .B1(n23725), .B2(n24327), .O(
        n23728) );
  OAI22S U28962 ( .A1(n30456), .A2(n24319), .B1(n24272), .B2(n24270), .O(
        n23727) );
  AO12 U28963 ( .B1(n23729), .B2(n23728), .A1(n23727), .O(n23734) );
  NR2 U28964 ( .I1(mem_data_out_reg_shift_1[22]), .I2(n23730), .O(n23732) );
  NR2 U28965 ( .I1(mem_data_out_reg_shift_1[23]), .I2(n24340), .O(n23731) );
  NR2 U28966 ( .I1(n23732), .I2(n23731), .O(n23733) );
  AOI22H U28967 ( .A1(mem_data_out_reg_shift_1[23]), .A2(n23954), .B1(n23734), 
        .B2(n23733), .O(n23737) );
  NR2F U28968 ( .I1(n23737), .I2(n23735), .O(n24604) );
  NR2T U28969 ( .I1(n23736), .I2(n24604), .O(n24616) );
  OR2T U28970 ( .I1(n24325), .I2(n24616), .O(n23963) );
  NR2F U28971 ( .I1(n23737), .I2(n23736), .O(n24263) );
  NR2T U28972 ( .I1(n24604), .I2(n23738), .O(n24614) );
  ND2S U28973 ( .I1(n23961), .I2(mem_data_out_reg_shift_1[19]), .O(n23739) );
  OAI12HS U28974 ( .B1(n23963), .B2(n24281), .A1(n23739), .O(n23741) );
  INV1S U28975 ( .I(n24285), .O(n24540) );
  OR2T U28976 ( .I1(n24604), .I2(n24262), .O(n23960) );
  NR2 U28977 ( .I1(n24540), .I2(n23960), .O(n23740) );
  NR2 U28978 ( .I1(n23741), .I2(n23740), .O(n24181) );
  INV1S U28979 ( .I(n24181), .O(n24460) );
  OR2T U28980 ( .I1(n23863), .I2(n30241), .O(n24918) );
  ND2S U28981 ( .I1(n24918), .I2(mem_data_out_reg_shift_0[19]), .O(n23742) );
  AOI22S U28982 ( .A1(n23984), .A2(mem_data_out_reg_shift_1[27]), .B1(n23782), 
        .B2(mem_data_out_reg_shift_0[27]), .O(n23745) );
  ND2S U28983 ( .I1(n23783), .I2(mem_data_out_reg_shift_0[19]), .O(n23744) );
  ND2S U28984 ( .I1(n23784), .I2(mem_data_out_reg_shift_1[19]), .O(n23743) );
  ND3P U28985 ( .I1(n23745), .I2(n23744), .I3(n23743), .O(n24541) );
  INV2 U28986 ( .I(n24541), .O(n24280) );
  ND2S U28987 ( .I1(n24918), .I2(mem_data_out_reg_shift_0[18]), .O(n23746) );
  AOI22S U28988 ( .A1(n23784), .A2(mem_data_out_reg_shift_1[18]), .B1(n23782), 
        .B2(mem_data_out_reg_shift_0[26]), .O(n23749) );
  ND2S U28989 ( .I1(n23783), .I2(mem_data_out_reg_shift_0[18]), .O(n23748) );
  ND2S U28990 ( .I1(n23984), .I2(mem_data_out_reg_shift_1[26]), .O(n23747) );
  INV1S U28991 ( .I(n24546), .O(n24289) );
  NR2 U28992 ( .I1(n24547), .I2(n24289), .O(n23750) );
  NR2 U28993 ( .I1(n23763), .I2(n23750), .O(n23766) );
  ND2S U28994 ( .I1(n24918), .I2(mem_data_out_reg_shift_0[17]), .O(n23751) );
  AOI22S U28995 ( .A1(n23784), .A2(mem_data_out_reg_shift_1[17]), .B1(n23782), 
        .B2(mem_data_out_reg_shift_0[25]), .O(n23754) );
  ND2S U28996 ( .I1(n23783), .I2(mem_data_out_reg_shift_0[17]), .O(n23753) );
  ND2S U28997 ( .I1(n23984), .I2(mem_data_out_reg_shift_1[25]), .O(n23752) );
  INV2 U28998 ( .I(n24557), .O(n24299) );
  NR2 U28999 ( .I1(n24556), .I2(n24299), .O(n23760) );
  INV1S U29000 ( .I(mem_data_out_reg_shift_1[16]), .O(n24301) );
  ND2S U29001 ( .I1(n24918), .I2(mem_data_out_reg_shift_0[16]), .O(n23755) );
  OAI12HS U29002 ( .B1(n23781), .B2(n24301), .A1(n23755), .O(n24762) );
  ND2S U29003 ( .I1(n23783), .I2(mem_data_out_reg_shift_0[16]), .O(n23758) );
  AOI22S U29004 ( .A1(n23784), .A2(mem_data_out_reg_shift_1[16]), .B1(n23984), 
        .B2(mem_data_out_reg_shift_1[24]), .O(n23757) );
  ND2S U29005 ( .I1(n23782), .I2(mem_data_out_reg_shift_0[24]), .O(n23756) );
  ND2S U29006 ( .I1(n24299), .I2(n24556), .O(n23759) );
  OAI12HS U29007 ( .B1(n23760), .B2(n15981), .A1(n23759), .O(n23765) );
  ND2S U29008 ( .I1(n24289), .I2(n24547), .O(n23762) );
  ND2S U29009 ( .I1(n24280), .I2(n24542), .O(n23761) );
  OAI12HS U29010 ( .B1(n23763), .B2(n23762), .A1(n23761), .O(n23764) );
  ND2S U29011 ( .I1(n24918), .I2(mem_data_out_reg_shift_0[23]), .O(n23767) );
  OAI12H U29012 ( .B1(n23781), .B2(n24341), .A1(n23767), .O(n24600) );
  ND2S U29013 ( .I1(n23783), .I2(mem_data_out_reg_shift_0[23]), .O(n23770) );
  AOI22S U29014 ( .A1(n23784), .A2(mem_data_out_reg_shift_1[23]), .B1(n23984), 
        .B2(mem_data_out_reg_shift_1[31]), .O(n23769) );
  ND2S U29015 ( .I1(n23782), .I2(mem_data_out_reg_shift_0[31]), .O(n23768) );
  ND2S U29016 ( .I1(n24918), .I2(mem_data_out_reg_shift_0[22]), .O(n23771) );
  AOI22S U29017 ( .A1(n23984), .A2(mem_data_out_reg_shift_1[30]), .B1(n23782), 
        .B2(mem_data_out_reg_shift_0[30]), .O(n23774) );
  ND2S U29018 ( .I1(n23783), .I2(mem_data_out_reg_shift_0[22]), .O(n23773) );
  ND2S U29019 ( .I1(n23784), .I2(mem_data_out_reg_shift_1[22]), .O(n23772) );
  NR2 U29020 ( .I1(n24609), .I2(n24276), .O(n23775) );
  ND2S U29021 ( .I1(n24918), .I2(mem_data_out_reg_shift_0[21]), .O(n23776) );
  AOI22S U29022 ( .A1(n23784), .A2(mem_data_out_reg_shift_1[21]), .B1(n23782), 
        .B2(mem_data_out_reg_shift_0[29]), .O(n23779) );
  ND2S U29023 ( .I1(n23783), .I2(mem_data_out_reg_shift_0[21]), .O(n23778) );
  ND2S U29024 ( .I1(n23984), .I2(mem_data_out_reg_shift_1[29]), .O(n23777) );
  ND3P U29025 ( .I1(n23779), .I2(n23778), .I3(n23777), .O(n24588) );
  INV1S U29026 ( .I(n24588), .O(n24315) );
  AOI22S U29027 ( .A1(n23984), .A2(mem_data_out_reg_shift_1[28]), .B1(n23782), 
        .B2(mem_data_out_reg_shift_0[28]), .O(n23787) );
  ND2S U29028 ( .I1(n23783), .I2(mem_data_out_reg_shift_0[20]), .O(n23786) );
  ND2S U29029 ( .I1(n23784), .I2(mem_data_out_reg_shift_1[20]), .O(n23785) );
  INV1 U29030 ( .I(n24578), .O(n24323) );
  NR2 U29031 ( .I1(n24579), .I2(n24323), .O(n23788) );
  NR2 U29032 ( .I1(n23792), .I2(n23788), .O(n23789) );
  ND2S U29033 ( .I1(n24323), .I2(n24579), .O(n23791) );
  OAI12HS U29034 ( .B1(n23792), .B2(n23791), .A1(n23790), .O(n23797) );
  ND2S U29035 ( .I1(n24276), .I2(n24609), .O(n23794) );
  ND2S U29036 ( .I1(n23950), .I2(n24600), .O(n23793) );
  ND2S U29037 ( .I1(n30241), .I2(mem_data_out_reg_shift_0[19]), .O(n23806) );
  MOAI1S U29038 ( .A1(n24919), .A2(n23802), .B1(medfilt_state[3]), .B2(
        mem_data_out_reg_shift_1[19]), .O(n23803) );
  INV1S U29039 ( .I(n23803), .O(n23805) );
  ND2S U29040 ( .I1(n23863), .I2(mem_data_out_reg_shift_0[11]), .O(n23804) );
  ND3 U29041 ( .I1(n23806), .I2(n23805), .I3(n23804), .O(n24277) );
  NR2 U29042 ( .I1(n24545), .I2(n24541), .O(n23822) );
  ND2S U29043 ( .I1(n30241), .I2(mem_data_out_reg_shift_0[18]), .O(n23811) );
  MOAI1S U29044 ( .A1(n24919), .A2(n23807), .B1(medfilt_state[3]), .B2(
        mem_data_out_reg_shift_1[18]), .O(n23808) );
  INV1S U29045 ( .I(n23808), .O(n23810) );
  ND2S U29046 ( .I1(n23863), .I2(mem_data_out_reg_shift_0[10]), .O(n23809) );
  NR2 U29047 ( .I1(n24550), .I2(n24546), .O(n23812) );
  NR2 U29048 ( .I1(n23822), .I2(n23812), .O(n23825) );
  ND2S U29049 ( .I1(n30241), .I2(mem_data_out_reg_shift_0[17]), .O(n23817) );
  MOAI1S U29050 ( .A1(n24919), .A2(n23813), .B1(medfilt_state[3]), .B2(
        mem_data_out_reg_shift_1[17]), .O(n23814) );
  INV1S U29051 ( .I(n23814), .O(n23816) );
  ND2S U29052 ( .I1(n23863), .I2(mem_data_out_reg_shift_0[9]), .O(n23815) );
  NR2 U29053 ( .I1(n24560), .I2(n24856), .O(n23819) );
  ND2S U29054 ( .I1(n24856), .I2(n24560), .O(n23818) );
  OAI12HS U29055 ( .B1(n23819), .B2(n24299), .A1(n23818), .O(n23824) );
  ND2S U29056 ( .I1(n24546), .I2(n24550), .O(n23821) );
  ND2S U29057 ( .I1(n24541), .I2(n24545), .O(n23820) );
  OAI12HS U29058 ( .B1(n23822), .B2(n23821), .A1(n23820), .O(n23823) );
  AOI12HS U29059 ( .B1(n23825), .B2(n23824), .A1(n23823), .O(n23860) );
  ND2S U29060 ( .I1(n30241), .I2(mem_data_out_reg_shift_0[21]), .O(n23830) );
  MOAI1S U29061 ( .A1(n24919), .A2(n23826), .B1(mem_data_out_reg_shift_1[21]), 
        .B2(medfilt_state[3]), .O(n23827) );
  INV1S U29062 ( .I(n23827), .O(n23829) );
  ND2S U29063 ( .I1(n23863), .I2(mem_data_out_reg_shift_0[13]), .O(n23828) );
  NR2 U29064 ( .I1(n24592), .I2(n24588), .O(n23851) );
  ND2S U29065 ( .I1(n30241), .I2(mem_data_out_reg_shift_0[20]), .O(n23835) );
  MOAI1S U29066 ( .A1(n24919), .A2(n23831), .B1(medfilt_state[3]), .B2(
        mem_data_out_reg_shift_1[20]), .O(n23832) );
  INV1S U29067 ( .I(n23832), .O(n23834) );
  ND2S U29068 ( .I1(n23863), .I2(mem_data_out_reg_shift_0[12]), .O(n23833) );
  NR2 U29069 ( .I1(n24582), .I2(n24578), .O(n23836) );
  NR2 U29070 ( .I1(n23851), .I2(n23836), .O(n23848) );
  ND2S U29071 ( .I1(n30241), .I2(mem_data_out_reg_shift_0[22]), .O(n23841) );
  MOAI1S U29072 ( .A1(n24919), .A2(n23837), .B1(mem_data_out_reg_shift_1[22]), 
        .B2(medfilt_state[3]), .O(n23838) );
  INV1S U29073 ( .I(n23838), .O(n23840) );
  ND2S U29074 ( .I1(n23863), .I2(mem_data_out_reg_shift_0[14]), .O(n23839) );
  NR2 U29075 ( .I1(n24613), .I2(n24607), .O(n23847) );
  ND2S U29076 ( .I1(n30241), .I2(mem_data_out_reg_shift_0[23]), .O(n23846) );
  MOAI1S U29077 ( .A1(n24919), .A2(n23842), .B1(mem_data_out_reg_shift_1[23]), 
        .B2(medfilt_state[3]), .O(n23843) );
  INV1S U29078 ( .I(n23843), .O(n23845) );
  ND2S U29079 ( .I1(n23863), .I2(mem_data_out_reg_shift_0[15]), .O(n23844) );
  ND3 U29080 ( .I1(n23846), .I2(n23845), .I3(n23844), .O(n24598) );
  NR2 U29081 ( .I1(n23951), .I2(n24599), .O(n23854) );
  ND2S U29082 ( .I1(n24588), .I2(n24592), .O(n23849) );
  OAI12HS U29083 ( .B1(n23851), .B2(n23850), .A1(n23849), .O(n23856) );
  ND2S U29084 ( .I1(n24607), .I2(n24613), .O(n23853) );
  ND2S U29085 ( .I1(n24599), .I2(n23951), .O(n23852) );
  OAI12HS U29086 ( .B1(n23854), .B2(n23853), .A1(n23852), .O(n23855) );
  AOI12HS U29087 ( .B1(n23857), .B2(n23856), .A1(n23855), .O(n23858) );
  NR2 U29088 ( .I1(n24545), .I2(n24542), .O(n23872) );
  NR2 U29089 ( .I1(n24550), .I2(n24547), .O(n23861) );
  NR2 U29090 ( .I1(n23872), .I2(n23861), .O(n23875) );
  ND2S U29091 ( .I1(n30241), .I2(mem_data_out_reg_shift_0[16]), .O(n23866) );
  INV1S U29092 ( .I(mem_data_out_reg_shift_1[8]), .O(n23904) );
  MOAI1S U29093 ( .A1(n24919), .A2(n23904), .B1(medfilt_state[3]), .B2(
        mem_data_out_reg_shift_1[16]), .O(n23862) );
  INV1S U29094 ( .I(n23862), .O(n23865) );
  ND2S U29095 ( .I1(n23863), .I2(mem_data_out_reg_shift_0[8]), .O(n23864) );
  ND3S U29096 ( .I1(n23866), .I2(n23865), .I3(n23864), .O(n24760) );
  INV1S U29097 ( .I(n24760), .O(n24861) );
  NR2 U29098 ( .I1(n24861), .I2(n24560), .O(n23869) );
  INV1S U29099 ( .I(n24556), .O(n23868) );
  ND2S U29100 ( .I1(n24560), .I2(n24861), .O(n23867) );
  OAI12HS U29101 ( .B1(n23869), .B2(n23868), .A1(n23867), .O(n23874) );
  ND2S U29102 ( .I1(n24547), .I2(n24550), .O(n23871) );
  ND2S U29103 ( .I1(n24542), .I2(n24545), .O(n23870) );
  OAI12HS U29104 ( .B1(n23872), .B2(n23871), .A1(n23870), .O(n23873) );
  NR2 U29105 ( .I1(n24582), .I2(n24579), .O(n23876) );
  NR2 U29106 ( .I1(n23881), .I2(n23876), .O(n23878) );
  NR2 U29107 ( .I1(n24613), .I2(n24609), .O(n23877) );
  NR2 U29108 ( .I1(n23884), .I2(n23877), .O(n23887) );
  ND2S U29109 ( .I1(n24579), .I2(n24582), .O(n23880) );
  OAI12HS U29110 ( .B1(n23881), .B2(n23880), .A1(n23879), .O(n23886) );
  ND2S U29111 ( .I1(n24609), .I2(n24613), .O(n23883) );
  ND2S U29112 ( .I1(n24600), .I2(n23951), .O(n23882) );
  OAI12HS U29113 ( .B1(n23884), .B2(n23883), .A1(n23882), .O(n23885) );
  NR2P U29114 ( .I1(n24427), .I2(n24862), .O(n23937) );
  ND2S U29115 ( .I1(n23937), .I2(n24542), .O(n23894) );
  NR2P U29116 ( .I1(n24430), .I2(n24862), .O(n23939) );
  ND2S U29117 ( .I1(n23939), .I2(n24541), .O(n23893) );
  AOI22S U29118 ( .A1(n23946), .A2(n24541), .B1(n23938), .B2(n24542), .O(
        n23892) );
  ND3S U29119 ( .I1(n23894), .I2(n23893), .I3(n23892), .O(n23898) );
  NR2F U29120 ( .I1(n23896), .I2(n24430), .O(n24763) );
  NR2T U29121 ( .I1(n24764), .I2(n24763), .O(n24761) );
  NR2 U29122 ( .I1(n24545), .I2(n24434), .O(n23897) );
  NR2T U29123 ( .I1(n23898), .I2(n23897), .O(n24458) );
  ND2S U29124 ( .I1(n23937), .I2(n24556), .O(n23901) );
  ND2S U29125 ( .I1(n23939), .I2(n24557), .O(n23900) );
  AOI22S U29126 ( .A1(n23946), .A2(n24557), .B1(n23938), .B2(n24556), .O(
        n23899) );
  ND3S U29127 ( .I1(n23901), .I2(n23900), .I3(n23899), .O(n23903) );
  NR2 U29128 ( .I1(n24560), .I2(n24434), .O(n23902) );
  NR2 U29129 ( .I1(n23903), .I2(n23902), .O(n24226) );
  INV1S U29130 ( .I(n24226), .O(n24258) );
  INV1S U29131 ( .I(n23960), .O(n23907) );
  OAI22S U29132 ( .A1(n24301), .A2(n23906), .B1(n23905), .B2(n23904), .O(
        n24561) );
  ND2S U29133 ( .I1(n23907), .I2(n24561), .O(n23912) );
  ND2S U29134 ( .I1(n23961), .I2(mem_data_out_reg_shift_1[16]), .O(n23911) );
  INV1S U29135 ( .I(n23963), .O(n23909) );
  INV1S U29136 ( .I(n23908), .O(n24562) );
  ND2S U29137 ( .I1(n23909), .I2(n24562), .O(n23910) );
  ND3 U29138 ( .I1(n23912), .I2(n23911), .I3(n23910), .O(n24426) );
  INV1S U29139 ( .I(n24426), .O(n23917) );
  INV1S U29140 ( .I(n24267), .O(n24569) );
  NR2 U29141 ( .I1(n24569), .I2(n23960), .O(n23916) );
  ND2S U29142 ( .I1(n23961), .I2(mem_data_out_reg_shift_1[17]), .O(n23913) );
  OAI12HS U29143 ( .B1(n23963), .B2(n23914), .A1(n23913), .O(n23915) );
  NR2P U29144 ( .I1(n23916), .I2(n23915), .O(n24223) );
  MAO222 U29145 ( .A1(n24258), .B1(n23917), .C1(n24223), .O(n23927) );
  ND2S U29146 ( .I1(n23937), .I2(n24547), .O(n23920) );
  ND2S U29147 ( .I1(n23939), .I2(n24546), .O(n23919) );
  AOI22S U29148 ( .A1(n23946), .A2(n24546), .B1(n23938), .B2(n24547), .O(
        n23918) );
  ND3S U29149 ( .I1(n23920), .I2(n23919), .I3(n23918), .O(n23922) );
  NR2 U29150 ( .I1(n24550), .I2(n24434), .O(n23921) );
  NR2P U29151 ( .I1(n23922), .I2(n23921), .O(n24447) );
  INV1S U29152 ( .I(n24294), .O(n24554) );
  NR2 U29153 ( .I1(n24554), .I2(n23960), .O(n23925) );
  ND2S U29154 ( .I1(n23961), .I2(mem_data_out_reg_shift_1[18]), .O(n23923) );
  OAI12HS U29155 ( .B1(n23963), .B2(n24290), .A1(n23923), .O(n23924) );
  NR2 U29156 ( .I1(n23925), .I2(n23924), .O(n24180) );
  INV1 U29157 ( .I(n24180), .O(n24446) );
  NR2 U29158 ( .I1(n24447), .I2(n24446), .O(n23926) );
  MOAI1 U29159 ( .A1(n23927), .A2(n23926), .B1(n24447), .B2(n24446), .O(n23936) );
  ND2S U29160 ( .I1(n23937), .I2(n24579), .O(n23930) );
  ND2S U29161 ( .I1(n23939), .I2(n24578), .O(n23929) );
  AOI22S U29162 ( .A1(n23946), .A2(n24578), .B1(n23938), .B2(n24579), .O(
        n23928) );
  ND3S U29163 ( .I1(n23930), .I2(n23929), .I3(n23928), .O(n23932) );
  NR2 U29164 ( .I1(n24582), .I2(n24434), .O(n23931) );
  NR2 U29165 ( .I1(n23932), .I2(n23931), .O(n24236) );
  INV1S U29166 ( .I(n24236), .O(n24503) );
  INV1S U29167 ( .I(n24330), .O(n24587) );
  NR2 U29168 ( .I1(n24587), .I2(n23960), .O(n23935) );
  ND2S U29169 ( .I1(n23961), .I2(mem_data_out_reg_shift_1[20]), .O(n23933) );
  OAI12HS U29170 ( .B1(n23963), .B2(n24324), .A1(n23933), .O(n23934) );
  NR2P U29171 ( .I1(n23935), .I2(n23934), .O(n24501) );
  ND2S U29172 ( .I1(n24503), .I2(n24501), .O(n23972) );
  OAI112HS U29173 ( .C1(n24460), .C2(n24458), .A1(n23936), .B1(n23972), .O(
        n23983) );
  OR2 U29174 ( .I1(n24613), .I2(n24434), .O(n23942) );
  ND2S U29175 ( .I1(n23966), .I2(n24609), .O(n23941) );
  ND2S U29176 ( .I1(n23967), .I2(n24607), .O(n23940) );
  INV1S U29177 ( .I(n24272), .O(n24619) );
  NR2 U29178 ( .I1(n24619), .I2(n23960), .O(n23945) );
  ND2S U29179 ( .I1(n23961), .I2(mem_data_out_reg_shift_1[22]), .O(n23943) );
  OAI12HS U29180 ( .B1(n23963), .B2(n24268), .A1(n23943), .O(n23944) );
  NR2P U29181 ( .I1(n23945), .I2(n23944), .O(n24478) );
  NR2 U29182 ( .I1(n24480), .I2(n24478), .O(n23959) );
  ND2S U29183 ( .I1(n23946), .I2(n24599), .O(n23948) );
  INV1S U29184 ( .I(n24600), .O(n23947) );
  AOI22S U29185 ( .A1(n23950), .A2(n23949), .B1(n23948), .B2(n23947), .O(
        n23953) );
  NR2 U29186 ( .I1(n23951), .I2(n24434), .O(n23952) );
  NR2 U29187 ( .I1(n23953), .I2(n23952), .O(n24245) );
  INV1S U29188 ( .I(n24245), .O(n24489) );
  ND2S U29189 ( .I1(n23961), .I2(mem_data_out_reg_shift_1[23]), .O(n23955) );
  OAI12HS U29190 ( .B1(n23963), .B2(n23956), .A1(n23955), .O(n23957) );
  NR2P U29191 ( .I1(n23958), .I2(n23957), .O(n24487) );
  NR2 U29192 ( .I1(n24489), .I2(n24487), .O(n23978) );
  NR2 U29193 ( .I1(n23959), .I2(n23978), .O(n23982) );
  INV1S U29194 ( .I(n24319), .O(n24596) );
  NR2 U29195 ( .I1(n24596), .I2(n23960), .O(n23965) );
  ND2S U29196 ( .I1(n23961), .I2(mem_data_out_reg_shift_1[21]), .O(n23962) );
  OAI12HS U29197 ( .B1(n23963), .B2(n24316), .A1(n23962), .O(n23964) );
  NR2P U29198 ( .I1(n23965), .I2(n23964), .O(n24515) );
  OR2 U29199 ( .I1(n24592), .I2(n24434), .O(n23970) );
  ND2S U29200 ( .I1(n23967), .I2(n24588), .O(n23968) );
  ND3 U29201 ( .I1(n23970), .I2(n23969), .I3(n23968), .O(n24518) );
  OAI22S U29202 ( .A1(n24501), .A2(n24503), .B1(n24515), .B2(n24518), .O(
        n23971) );
  AOI13HS U29203 ( .B1(n24458), .B2(n23972), .B3(n24460), .A1(n23971), .O(
        n23981) );
  INV1S U29204 ( .I(n24480), .O(n23974) );
  INV1S U29205 ( .I(n24518), .O(n23973) );
  NR2 U29206 ( .I1(n23974), .I2(n23973), .O(n23977) );
  ND2S U29207 ( .I1(n24515), .I2(n24518), .O(n23975) );
  ND2S U29208 ( .I1(n23975), .I2(n23974), .O(n23976) );
  AOI22S U29209 ( .A1(n23977), .A2(n24515), .B1(n23976), .B2(n24478), .O(
        n23979) );
  MOAI1 U29210 ( .A1(n23979), .A2(n23978), .B1(n24487), .B2(n24489), .O(n23980) );
  AOI13H U29211 ( .B1(n23983), .B2(n23982), .B3(n23981), .A1(n23980), .O(
        n24253) );
  INV1S U29212 ( .I(mem_data_out_reg_shift_2[27]), .O(n23985) );
  NR2F U29213 ( .I1(n24928), .I2(n23984), .O(n24041) );
  NR2 U29214 ( .I1(n23985), .I2(n24041), .O(n23991) );
  OR2P U29215 ( .I1(n23987), .I2(n23986), .O(n24043) );
  ND2S U29216 ( .I1(n24043), .I2(mem_data_out_reg_shift_2[19]), .O(n23989) );
  OR2P U29217 ( .I1(n24100), .I2(n24909), .O(n24044) );
  ND2S U29218 ( .I1(n24044), .I2(mem_data_out_reg_shift_1[27]), .O(n23988) );
  OAI112HS U29219 ( .C1(n24283), .C2(n24047), .A1(n23989), .B1(n23988), .O(
        n23990) );
  INV2 U29220 ( .I(n24041), .O(n23992) );
  NR2F U29221 ( .I1(n24043), .I2(n23992), .O(n24052) );
  INV1S U29222 ( .I(mem_data_out_reg_shift_2[16]), .O(n23994) );
  INV1 U29223 ( .I(n23993), .O(n23996) );
  OR2T U29224 ( .I1(n23996), .I2(n24909), .O(n24114) );
  OR2P U29225 ( .I1(n24100), .I2(n24114), .O(n24050) );
  MOAI1H U29226 ( .A1(n24052), .A2(n23994), .B1(mem_data_out_reg_shift_1[16]), 
        .B2(n24050), .O(n24354) );
  INV2 U29227 ( .I(n24354), .O(n24652) );
  INV1S U29228 ( .I(mem_data_out_reg_shift_2[24]), .O(n23995) );
  AOI22S U29229 ( .A1(n23996), .A2(mem_data_out_reg_shift_1[16]), .B1(n24044), 
        .B2(mem_data_out_reg_shift_1[24]), .O(n23998) );
  ND2S U29230 ( .I1(n24043), .I2(mem_data_out_reg_shift_2[16]), .O(n23997) );
  ND3 U29231 ( .I1(n23999), .I2(n23998), .I3(n23997), .O(n24353) );
  INV1S U29232 ( .I(mem_data_out_reg_shift_2[25]), .O(n24000) );
  NR2 U29233 ( .I1(n24000), .I2(n24041), .O(n24004) );
  ND2S U29234 ( .I1(n24044), .I2(mem_data_out_reg_shift_1[25]), .O(n24002) );
  ND2S U29235 ( .I1(n24043), .I2(mem_data_out_reg_shift_2[17]), .O(n24001) );
  OAI112HS U29236 ( .C1(n24265), .C2(n24047), .A1(n24002), .B1(n24001), .O(
        n24003) );
  NR2T U29237 ( .I1(n24004), .I2(n24003), .O(n24660) );
  INV1S U29238 ( .I(mem_data_out_reg_shift_2[17]), .O(n24005) );
  MOAI1H U29239 ( .A1(n24052), .A2(n24005), .B1(mem_data_out_reg_shift_1[17]), 
        .B2(n24050), .O(n24658) );
  NR2 U29240 ( .I1(n24660), .I2(n24658), .O(n24007) );
  ND2S U29241 ( .I1(n24658), .I2(n24660), .O(n24006) );
  INV1S U29242 ( .I(mem_data_out_reg_shift_2[19]), .O(n24008) );
  MOAI1H U29243 ( .A1(n24052), .A2(n24008), .B1(mem_data_out_reg_shift_1[19]), 
        .B2(n24050), .O(n24644) );
  NR2 U29244 ( .I1(n24646), .I2(n24644), .O(n24018) );
  INV1S U29245 ( .I(mem_data_out_reg_shift_2[26]), .O(n24009) );
  NR2 U29246 ( .I1(n24009), .I2(n24041), .O(n24013) );
  ND2S U29247 ( .I1(n24043), .I2(mem_data_out_reg_shift_2[18]), .O(n24011) );
  ND2S U29248 ( .I1(n24044), .I2(mem_data_out_reg_shift_1[26]), .O(n24010) );
  OAI112HS U29249 ( .C1(n24292), .C2(n24047), .A1(n24011), .B1(n24010), .O(
        n24012) );
  INV1S U29250 ( .I(mem_data_out_reg_shift_2[18]), .O(n24014) );
  MOAI1H U29251 ( .A1(n24052), .A2(n24014), .B1(mem_data_out_reg_shift_1[18]), 
        .B2(n24050), .O(n24636) );
  NR2 U29252 ( .I1(n24638), .I2(n24636), .O(n24015) );
  NR2 U29253 ( .I1(n24018), .I2(n24015), .O(n24020) );
  ND2S U29254 ( .I1(n24636), .I2(n24638), .O(n24017) );
  ND2S U29255 ( .I1(n24644), .I2(n24646), .O(n24016) );
  OAI12HS U29256 ( .B1(n24018), .B2(n24017), .A1(n24016), .O(n24019) );
  INV1S U29257 ( .I(mem_data_out_reg_shift_2[28]), .O(n24022) );
  NR2 U29258 ( .I1(n24022), .I2(n24041), .O(n24026) );
  ND2S U29259 ( .I1(n24043), .I2(mem_data_out_reg_shift_2[20]), .O(n24024) );
  ND2S U29260 ( .I1(n24044), .I2(mem_data_out_reg_shift_1[28]), .O(n24023) );
  OAI112HS U29261 ( .C1(n24327), .C2(n24047), .A1(n24024), .B1(n24023), .O(
        n24025) );
  NR2P U29262 ( .I1(n24026), .I2(n24025), .O(n24688) );
  INV1S U29263 ( .I(mem_data_out_reg_shift_2[20]), .O(n24027) );
  MOAI1H U29264 ( .A1(n24052), .A2(n24027), .B1(mem_data_out_reg_shift_1[20]), 
        .B2(n24050), .O(n24686) );
  NR2 U29265 ( .I1(n24688), .I2(n24686), .O(n24034) );
  INV1S U29266 ( .I(mem_data_out_reg_shift_2[29]), .O(n24028) );
  NR2 U29267 ( .I1(n24028), .I2(n24041), .O(n24032) );
  ND2S U29268 ( .I1(n24043), .I2(mem_data_out_reg_shift_2[21]), .O(n24030) );
  ND2S U29269 ( .I1(n24044), .I2(mem_data_out_reg_shift_1[29]), .O(n24029) );
  OAI112HS U29270 ( .C1(n30456), .C2(n24047), .A1(n24030), .B1(n24029), .O(
        n24031) );
  NR2P U29271 ( .I1(n24032), .I2(n24031), .O(n24696) );
  INV1S U29272 ( .I(mem_data_out_reg_shift_2[21]), .O(n24033) );
  MOAI1H U29273 ( .A1(n24052), .A2(n24033), .B1(mem_data_out_reg_shift_1[21]), 
        .B2(n24050), .O(n24378) );
  NR2 U29274 ( .I1(n24696), .I2(n24378), .O(n24057) );
  NR2 U29275 ( .I1(n24034), .I2(n24057), .O(n24054) );
  INV1S U29276 ( .I(mem_data_out_reg_shift_2[31]), .O(n24035) );
  NR2 U29277 ( .I1(n24035), .I2(n24041), .O(n24039) );
  ND2S U29278 ( .I1(n24043), .I2(mem_data_out_reg_shift_2[23]), .O(n24037) );
  ND2S U29279 ( .I1(n24044), .I2(mem_data_out_reg_shift_1[31]), .O(n24036) );
  OAI112HS U29280 ( .C1(n24047), .C2(n24341), .A1(n24037), .B1(n24036), .O(
        n24038) );
  INV1S U29281 ( .I(mem_data_out_reg_shift_2[23]), .O(n24040) );
  MOAI1H U29282 ( .A1(n24052), .A2(n24040), .B1(mem_data_out_reg_shift_1[23]), 
        .B2(n24050), .O(n24676) );
  INV1S U29283 ( .I(mem_data_out_reg_shift_2[30]), .O(n24042) );
  NR2 U29284 ( .I1(n24042), .I2(n24041), .O(n24049) );
  ND2S U29285 ( .I1(n24043), .I2(mem_data_out_reg_shift_2[22]), .O(n24046) );
  ND2S U29286 ( .I1(n24044), .I2(mem_data_out_reg_shift_1[30]), .O(n24045) );
  OAI112HS U29287 ( .C1(n24270), .C2(n24047), .A1(n24046), .B1(n24045), .O(
        n24048) );
  NR2P U29288 ( .I1(n24049), .I2(n24048), .O(n24680) );
  INV1S U29289 ( .I(mem_data_out_reg_shift_2[22]), .O(n24051) );
  NR2 U29290 ( .I1(n24680), .I2(n24345), .O(n24053) );
  ND2 U29291 ( .I1(n24054), .I2(n24063), .O(n24065) );
  ND2S U29292 ( .I1(n24686), .I2(n24688), .O(n24056) );
  ND2S U29293 ( .I1(n24378), .I2(n24696), .O(n24055) );
  OAI12HS U29294 ( .B1(n24057), .B2(n24056), .A1(n24055), .O(n24062) );
  ND2S U29295 ( .I1(n24345), .I2(n24680), .O(n24059) );
  ND2S U29296 ( .I1(n24676), .I2(n24674), .O(n24058) );
  OAI12HS U29297 ( .B1(n24060), .B2(n24059), .A1(n24058), .O(n24061) );
  INV1S U29298 ( .I(mem_data_out_reg_shift_2[11]), .O(n24070) );
  ND2P U29299 ( .I1(n24068), .I2(n24067), .O(n24927) );
  NR2F U29300 ( .I1(n24069), .I2(n24927), .O(n24119) );
  OR2 U29301 ( .I1(n24070), .I2(n24119), .O(n24073) );
  AOI22S U29302 ( .A1(n24100), .A2(mem_data_out_reg_shift_1[19]), .B1(n24115), 
        .B2(mem_data_out_reg_shift_2[19]), .O(n24072) );
  ND2S U29303 ( .I1(n24114), .I2(mem_data_out_reg_shift_1[11]), .O(n24071) );
  ND3P U29304 ( .I1(n24073), .I2(n24072), .I3(n24071), .O(n24647) );
  INV1S U29305 ( .I(n24647), .O(n24092) );
  NR2 U29306 ( .I1(n24092), .I2(n24644), .O(n24095) );
  INV1S U29307 ( .I(mem_data_out_reg_shift_2[10]), .O(n24074) );
  OR2 U29308 ( .I1(n24074), .I2(n24119), .O(n24077) );
  AOI22S U29309 ( .A1(n24100), .A2(mem_data_out_reg_shift_1[18]), .B1(n24114), 
        .B2(mem_data_out_reg_shift_1[10]), .O(n24076) );
  ND2S U29310 ( .I1(n24115), .I2(mem_data_out_reg_shift_2[18]), .O(n24075) );
  ND3P U29311 ( .I1(n24077), .I2(n24076), .I3(n24075), .O(n24640) );
  INV1S U29312 ( .I(n24640), .O(n24091) );
  NR2 U29313 ( .I1(n24091), .I2(n24636), .O(n24078) );
  NR2 U29314 ( .I1(n24095), .I2(n24078), .O(n24098) );
  INV1S U29315 ( .I(mem_data_out_reg_shift_2[9]), .O(n24079) );
  OR2 U29316 ( .I1(n24079), .I2(n24119), .O(n24082) );
  AOI22S U29317 ( .A1(n24100), .A2(mem_data_out_reg_shift_1[17]), .B1(n24114), 
        .B2(mem_data_out_reg_shift_1[9]), .O(n24081) );
  ND2S U29318 ( .I1(n24115), .I2(mem_data_out_reg_shift_2[17]), .O(n24080) );
  ND3P U29319 ( .I1(n24082), .I2(n24081), .I3(n24080), .O(n24661) );
  INV1S U29320 ( .I(n24661), .O(n24087) );
  NR2 U29321 ( .I1(n24087), .I2(n24658), .O(n24090) );
  INV1S U29322 ( .I(mem_data_out_reg_shift_2[8]), .O(n24083) );
  AOI22S U29323 ( .A1(n24100), .A2(mem_data_out_reg_shift_1[16]), .B1(n24114), 
        .B2(mem_data_out_reg_shift_1[8]), .O(n24085) );
  ND2S U29324 ( .I1(n24115), .I2(mem_data_out_reg_shift_2[16]), .O(n24084) );
  ND3P U29325 ( .I1(n24086), .I2(n24085), .I3(n24084), .O(n24654) );
  OR2 U29326 ( .I1(n24654), .I2(n24652), .O(n24089) );
  ND2S U29327 ( .I1(n24658), .I2(n24087), .O(n24088) );
  OAI12HS U29328 ( .B1(n24090), .B2(n24089), .A1(n24088), .O(n24097) );
  ND2S U29329 ( .I1(n24636), .I2(n24091), .O(n24094) );
  ND2S U29330 ( .I1(n24644), .I2(n24092), .O(n24093) );
  OAI12HS U29331 ( .B1(n24095), .B2(n24094), .A1(n24093), .O(n24096) );
  INV1S U29332 ( .I(mem_data_out_reg_shift_2[12]), .O(n24099) );
  OR2 U29333 ( .I1(n24099), .I2(n24119), .O(n24103) );
  AOI22S U29334 ( .A1(n24100), .A2(mem_data_out_reg_shift_1[20]), .B1(n24115), 
        .B2(mem_data_out_reg_shift_2[20]), .O(n24102) );
  ND2S U29335 ( .I1(n24114), .I2(mem_data_out_reg_shift_1[12]), .O(n24101) );
  ND3 U29336 ( .I1(n24103), .I2(n24102), .I3(n24101), .O(n24689) );
  INV1S U29337 ( .I(n24689), .O(n24125) );
  NR2 U29338 ( .I1(n24125), .I2(n24686), .O(n24109) );
  ND2S U29339 ( .I1(n24114), .I2(mem_data_out_reg_shift_1[13]), .O(n24105) );
  ND2S U29340 ( .I1(n24115), .I2(mem_data_out_reg_shift_2[21]), .O(n24104) );
  OAI112HS U29341 ( .C1(n24118), .C2(n30456), .A1(n24105), .B1(n24104), .O(
        n24108) );
  INV1S U29342 ( .I(mem_data_out_reg_shift_2[13]), .O(n24106) );
  NR2 U29343 ( .I1(n24106), .I2(n24119), .O(n24107) );
  NR2P U29344 ( .I1(n24108), .I2(n24107), .O(n24139) );
  NR2 U29345 ( .I1(n24139), .I2(n24378), .O(n24128) );
  NR2 U29346 ( .I1(n24109), .I2(n24128), .O(n24124) );
  ND2S U29347 ( .I1(n24114), .I2(mem_data_out_reg_shift_1[15]), .O(n24111) );
  ND2S U29348 ( .I1(n24115), .I2(mem_data_out_reg_shift_2[23]), .O(n24110) );
  OAI112HS U29349 ( .C1(n24118), .C2(n24341), .A1(n24111), .B1(n24110), .O(
        n24113) );
  NR2 U29350 ( .I1(n30455), .I2(n24119), .O(n24112) );
  NR2P U29351 ( .I1(n24113), .I2(n24112), .O(n24677) );
  NR2 U29352 ( .I1(n24677), .I2(n24676), .O(n24131) );
  ND2S U29353 ( .I1(n24114), .I2(mem_data_out_reg_shift_1[14]), .O(n24117) );
  ND2S U29354 ( .I1(n24115), .I2(mem_data_out_reg_shift_2[22]), .O(n24116) );
  OAI112HS U29355 ( .C1(n24118), .C2(n24270), .A1(n24117), .B1(n24116), .O(
        n24122) );
  INV1S U29356 ( .I(mem_data_out_reg_shift_2[14]), .O(n24120) );
  NR2 U29357 ( .I1(n24120), .I2(n24119), .O(n24121) );
  NR2 U29358 ( .I1(n24196), .I2(n24345), .O(n24123) );
  ND2 U29359 ( .I1(n24124), .I2(n24134), .O(n24136) );
  ND2S U29360 ( .I1(n24686), .I2(n24125), .O(n24127) );
  ND2S U29361 ( .I1(n24378), .I2(n24139), .O(n24126) );
  ND2S U29362 ( .I1(n24345), .I2(n24196), .O(n24130) );
  ND2S U29363 ( .I1(n24676), .I2(n24677), .O(n24129) );
  OAI12HS U29364 ( .B1(n24131), .B2(n24130), .A1(n24129), .O(n24132) );
  AOI12HS U29365 ( .B1(n24134), .B2(n24133), .A1(n24132), .O(n24135) );
  INV2 U29366 ( .I(n24203), .O(n24171) );
  INV1S U29367 ( .I(n24139), .O(n24697) );
  NR2 U29368 ( .I1(n24696), .I2(n24697), .O(n24138) );
  INV1S U29369 ( .I(n24680), .O(n24141) );
  INV1S U29370 ( .I(n24696), .O(n24140) );
  OAI22S U29371 ( .A1(n24196), .A2(n24141), .B1(n24140), .B2(n24139), .O(
        n24156) );
  NR2P U29372 ( .I1(n24647), .I2(n24646), .O(n24148) );
  NR2 U29373 ( .I1(n24640), .I2(n24638), .O(n24142) );
  INV1 U29374 ( .I(n24654), .O(n24143) );
  NR2P U29375 ( .I1(n24661), .I2(n24660), .O(n24145) );
  ND2 U29376 ( .I1(n24660), .I2(n24661), .O(n24144) );
  OAI12H U29377 ( .B1(n15988), .B2(n24145), .A1(n24144), .O(n24150) );
  ND2S U29378 ( .I1(n24638), .I2(n24640), .O(n24147) );
  ND2S U29379 ( .I1(n24646), .I2(n24647), .O(n24146) );
  OAI12HS U29380 ( .B1(n24148), .B2(n24147), .A1(n24146), .O(n24149) );
  NR2 U29381 ( .I1(n24689), .I2(n24688), .O(n24153) );
  ND2S U29382 ( .I1(n24688), .I2(n24689), .O(n24152) );
  OAI12H U29383 ( .B1(n24154), .B2(n24153), .A1(n24152), .O(n24155) );
  INV1S U29384 ( .I(n24677), .O(n24207) );
  MAO222P U29385 ( .A1(n24159), .B1(n24674), .C1(n24207), .O(n24168) );
  NR2F U29386 ( .I1(n24171), .I2(n24168), .O(n24639) );
  INV3 U29387 ( .I(n24169), .O(n24170) );
  ND2P U29388 ( .I1(n24168), .I2(n24170), .O(n24205) );
  OR2 U29389 ( .I1(n24646), .I2(n15922), .O(n24163) );
  OR2P U29390 ( .I1(n24170), .I2(n24203), .O(n24197) );
  ND2S U29391 ( .I1(n24188), .I2(n24644), .O(n24162) );
  ND2P U29392 ( .I1(n24205), .I2(n24197), .O(n24382) );
  ND2S U29393 ( .I1(n24208), .I2(n24647), .O(n24161) );
  ND3P U29394 ( .I1(n24163), .I2(n24162), .I3(n24161), .O(n24461) );
  NR2 U29395 ( .I1(n24461), .I2(n24181), .O(n24184) );
  ND2S U29396 ( .I1(n24208), .I2(n24640), .O(n24166) );
  ND2S U29397 ( .I1(n24188), .I2(n24636), .O(n24165) );
  OR2 U29398 ( .I1(n24638), .I2(n15922), .O(n24164) );
  ND3P U29399 ( .I1(n24166), .I2(n24165), .I3(n24164), .O(n24445) );
  NR2 U29400 ( .I1(n24180), .I2(n24445), .O(n24167) );
  NR2 U29401 ( .I1(n24184), .I2(n24167), .O(n24187) );
  ND2S U29402 ( .I1(n24208), .I2(n24654), .O(n24175) );
  OR2T U29403 ( .I1(n24170), .I2(n24639), .O(n24695) );
  OR2P U29404 ( .I1(n24169), .I2(n24168), .O(n24380) );
  ND3S U29405 ( .I1(n24695), .I2(n24380), .I3(n24353), .O(n24174) );
  OR2T U29406 ( .I1(n24169), .I2(n24639), .O(n24693) );
  NR2P U29407 ( .I1(n24171), .I2(n24170), .O(n24379) );
  INV1S U29408 ( .I(n24379), .O(n24172) );
  ND3P U29409 ( .I1(n24175), .I2(n24174), .I3(n24173), .O(n24425) );
  NR2 U29410 ( .I1(n24223), .I2(n24425), .O(n24179) );
  ND2S U29411 ( .I1(n24208), .I2(n24661), .O(n24177) );
  ND2S U29412 ( .I1(n24188), .I2(n24658), .O(n24176) );
  OAI112HS U29413 ( .C1(n15922), .C2(n24660), .A1(n24177), .B1(n24176), .O(
        n24254) );
  ND2S U29414 ( .I1(n24425), .I2(n24223), .O(n24178) );
  OAI12HS U29415 ( .B1(n24179), .B2(n24228), .A1(n24178), .O(n24186) );
  ND2S U29416 ( .I1(n24445), .I2(n24180), .O(n24183) );
  ND2S U29417 ( .I1(n24461), .I2(n24181), .O(n24182) );
  OAI12HS U29418 ( .B1(n24184), .B2(n24183), .A1(n24182), .O(n24185) );
  AOI12HS U29419 ( .B1(n24187), .B2(n24186), .A1(n24185), .O(n24222) );
  ND2S U29420 ( .I1(n24208), .I2(n24689), .O(n24191) );
  ND2S U29421 ( .I1(n24188), .I2(n24686), .O(n24190) );
  OR2 U29422 ( .I1(n24688), .I2(n15922), .O(n24189) );
  NR2 U29423 ( .I1(n24501), .I2(n24500), .O(n24195) );
  ND2S U29424 ( .I1(n24208), .I2(n24697), .O(n24194) );
  INV1S U29425 ( .I(n24378), .O(n24694) );
  AO12 U29426 ( .B1(n24198), .B2(n24197), .A1(n24694), .O(n24193) );
  OR2 U29427 ( .I1(n24696), .I2(n15922), .O(n24192) );
  ND3P U29428 ( .I1(n24194), .I2(n24193), .I3(n24192), .O(n24513) );
  NR2 U29429 ( .I1(n24515), .I2(n24513), .O(n24213) );
  NR2 U29430 ( .I1(n24195), .I2(n24213), .O(n24210) );
  INV1S U29431 ( .I(n24196), .O(n24681) );
  ND2S U29432 ( .I1(n24208), .I2(n24681), .O(n24202) );
  INV1S U29433 ( .I(n24345), .O(n24679) );
  NR2 U29434 ( .I1(n24478), .I2(n24477), .O(n24209) );
  ND2S U29435 ( .I1(n24203), .I2(n24674), .O(n24204) );
  MOAI1S U29436 ( .A1(n24205), .A2(n24674), .B1(n24676), .B2(n24204), .O(
        n24206) );
  NR2 U29437 ( .I1(n24487), .I2(n24486), .O(n24216) );
  NR2 U29438 ( .I1(n24209), .I2(n24216), .O(n24218) );
  ND2S U29439 ( .I1(n24210), .I2(n24218), .O(n24221) );
  ND2S U29440 ( .I1(n24500), .I2(n24501), .O(n24212) );
  ND2S U29441 ( .I1(n24513), .I2(n24515), .O(n24211) );
  OAI12HS U29442 ( .B1(n24213), .B2(n24212), .A1(n24211), .O(n24219) );
  ND2S U29443 ( .I1(n24477), .I2(n24478), .O(n24215) );
  ND2S U29444 ( .I1(n24486), .I2(n24487), .O(n24214) );
  OAI12HS U29445 ( .B1(n24216), .B2(n24215), .A1(n24214), .O(n24217) );
  AOI12HS U29446 ( .B1(n24219), .B2(n24218), .A1(n24217), .O(n24220) );
  OAI12HS U29447 ( .B1(n24222), .B2(n24221), .A1(n24220), .O(n24252) );
  NR2P U29448 ( .I1(n24253), .I2(n24252), .O(n24257) );
  OR2T U29449 ( .I1(n24257), .I2(n15987), .O(n24517) );
  INV1S U29450 ( .I(n24223), .O(n24224) );
  ND2S U29451 ( .I1(n24517), .I2(n24224), .O(n24261) );
  NR2P U29452 ( .I1(n24458), .I2(n24461), .O(n24232) );
  NR2 U29453 ( .I1(n24447), .I2(n24445), .O(n24225) );
  NR2 U29454 ( .I1(n24226), .I2(n24425), .O(n24229) );
  ND2S U29455 ( .I1(n24425), .I2(n24226), .O(n24227) );
  ND2S U29456 ( .I1(n24461), .I2(n24458), .O(n24230) );
  OAI12HS U29457 ( .B1(n24232), .B2(n24231), .A1(n24230), .O(n24233) );
  AOI12H U29458 ( .B1(n24235), .B2(n24234), .A1(n24233), .O(n24239) );
  NR2 U29459 ( .I1(n24236), .I2(n24500), .O(n24238) );
  ND2S U29460 ( .I1(n24500), .I2(n24236), .O(n24237) );
  OAI12H U29461 ( .B1(n24239), .B2(n24238), .A1(n24237), .O(n24241) );
  ND2S U29462 ( .I1(n24241), .I2(n24513), .O(n24240) );
  ND2P U29463 ( .I1(n24242), .I2(n15986), .O(n24244) );
  INV1S U29464 ( .I(n24477), .O(n24246) );
  ND2S U29465 ( .I1(n24486), .I2(n24245), .O(n24247) );
  OA12 U29466 ( .B1(n24246), .B2(n24480), .A1(n24247), .O(n24243) );
  ND2P U29467 ( .I1(n24244), .I2(n24243), .O(n24250) );
  ND3S U29468 ( .I1(n24247), .I2(n24246), .I3(n24480), .O(n24248) );
  ND3P U29469 ( .I1(n24250), .I2(n24249), .I3(n24248), .O(n24251) );
  MXL2H U29470 ( .A(n24253), .B(n24252), .S(n24251), .OB(n24255) );
  ND2S U29471 ( .I1(n24514), .I2(n24254), .O(n24260) );
  INV3 U29472 ( .I(n24255), .O(n24256) );
  NR2T U29473 ( .I1(n24257), .I2(n24256), .O(n24519) );
  ND2S U29474 ( .I1(n24519), .I2(n24258), .O(n24259) );
  BUF2 U29475 ( .I(n24262), .O(n24331) );
  ND2S U29476 ( .I1(n24325), .I2(n24566), .O(n24264) );
  OAI12HS U29477 ( .B1(n24328), .B2(n24265), .A1(n24264), .O(n24266) );
  AOI12HS U29478 ( .B1(n24331), .B2(n24267), .A1(n24266), .O(n24417) );
  INV1S U29479 ( .I(n24268), .O(n24615) );
  ND2S U29480 ( .I1(n24325), .I2(n24615), .O(n24269) );
  OAI12HS U29481 ( .B1(n24328), .B2(n24270), .A1(n24269), .O(n24271) );
  AOI12HS U29482 ( .B1(n24331), .B2(n24272), .A1(n24271), .O(n24471) );
  INV1 U29483 ( .I(n24764), .O(n24431) );
  ND2S U29484 ( .I1(n24761), .I2(n24273), .O(n24275) );
  ND2S U29485 ( .I1(n24763), .I2(n24609), .O(n24274) );
  OAI112HS U29486 ( .C1(n24276), .C2(n24431), .A1(n24275), .B1(n24274), .O(
        n24376) );
  ND2S U29487 ( .I1(n24763), .I2(n24542), .O(n24278) );
  OAI112HS U29488 ( .C1(n24280), .C2(n24431), .A1(n24279), .B1(n24278), .O(
        n24359) );
  INV1S U29489 ( .I(n24281), .O(n24537) );
  ND2S U29490 ( .I1(n24325), .I2(n24537), .O(n24282) );
  OAI12HS U29491 ( .B1(n24328), .B2(n24283), .A1(n24282), .O(n24284) );
  NR2 U29492 ( .I1(n24359), .I2(n24452), .O(n24308) );
  ND2S U29493 ( .I1(n24761), .I2(n24286), .O(n24288) );
  ND2S U29494 ( .I1(n24763), .I2(n24547), .O(n24287) );
  OAI112HS U29495 ( .C1(n24289), .C2(n24431), .A1(n24288), .B1(n24287), .O(
        n24361) );
  INV1S U29496 ( .I(n24290), .O(n24551) );
  ND2S U29497 ( .I1(n24325), .I2(n24551), .O(n24291) );
  OAI12HS U29498 ( .B1(n24328), .B2(n24292), .A1(n24291), .O(n24293) );
  NR2 U29499 ( .I1(n24361), .I2(n24439), .O(n24295) );
  NR2 U29500 ( .I1(n24308), .I2(n24295), .O(n24311) );
  ND2S U29501 ( .I1(n24761), .I2(n24296), .O(n24298) );
  ND2S U29502 ( .I1(n24763), .I2(n24556), .O(n24297) );
  OAI112HS U29503 ( .C1(n24299), .C2(n24431), .A1(n24298), .B1(n24297), .O(
        n24351) );
  ND2S U29504 ( .I1(n24325), .I2(n24562), .O(n24300) );
  OAI12HS U29505 ( .B1(n24328), .B2(n24301), .A1(n24300), .O(n24302) );
  AOI12HS U29506 ( .B1(n24331), .B2(n24561), .A1(n24302), .O(n24769) );
  NR2 U29507 ( .I1(n24351), .I2(n24769), .O(n24305) );
  INV1S U29508 ( .I(n24417), .O(n24304) );
  ND2S U29509 ( .I1(n24769), .I2(n24351), .O(n24303) );
  OAI12HS U29510 ( .B1(n24305), .B2(n24304), .A1(n24303), .O(n24310) );
  ND2S U29511 ( .I1(n24439), .I2(n24361), .O(n24307) );
  ND2S U29512 ( .I1(n24452), .I2(n24359), .O(n24306) );
  OAI12HS U29513 ( .B1(n24308), .B2(n24307), .A1(n24306), .O(n24309) );
  AOI12HS U29514 ( .B1(n24311), .B2(n24310), .A1(n24309), .O(n24338) );
  ND2S U29515 ( .I1(n24761), .I2(n24312), .O(n24314) );
  ND2S U29516 ( .I1(n24763), .I2(n24589), .O(n24313) );
  OAI112HS U29517 ( .C1(n24315), .C2(n24431), .A1(n24314), .B1(n24313), .O(
        n24375) );
  INV1S U29518 ( .I(n24316), .O(n24593) );
  ND2S U29519 ( .I1(n24325), .I2(n24593), .O(n24317) );
  OAI12HS U29520 ( .B1(n24328), .B2(n30456), .A1(n24317), .O(n24318) );
  NR2 U29521 ( .I1(n24375), .I2(n24507), .O(n24335) );
  ND2S U29522 ( .I1(n24761), .I2(n24320), .O(n24322) );
  ND2S U29523 ( .I1(n24763), .I2(n24579), .O(n24321) );
  OAI112HS U29524 ( .C1(n24323), .C2(n24431), .A1(n24322), .B1(n24321), .O(
        n24370) );
  INV1S U29525 ( .I(n24324), .O(n24584) );
  ND2S U29526 ( .I1(n24325), .I2(n24584), .O(n24326) );
  OAI12HS U29527 ( .B1(n24328), .B2(n24327), .A1(n24326), .O(n24329) );
  AOI12HS U29528 ( .B1(n24331), .B2(n24330), .A1(n24329), .O(n24494) );
  NR2 U29529 ( .I1(n24370), .I2(n24494), .O(n24332) );
  ND2S U29530 ( .I1(n24494), .I2(n24370), .O(n24334) );
  ND2S U29531 ( .I1(n24507), .I2(n24375), .O(n24333) );
  OAI12HS U29532 ( .B1(n24338), .B2(n24337), .A1(n24336), .O(n24343) );
  OR2S U29533 ( .I1(n24599), .I2(n24598), .O(n24339) );
  NR2 U29534 ( .I1(n24339), .I2(n24600), .O(n24485) );
  ND3S U29535 ( .I1(n24342), .I2(n24341), .I3(n24340), .O(n24400) );
  ND2S U29536 ( .I1(n24485), .I2(n24400), .O(n24348) );
  OAI112HS U29537 ( .C1(n24471), .C2(n24376), .A1(n24343), .B1(n24348), .O(
        n24389) );
  INV1S U29538 ( .I(n24485), .O(n24350) );
  INV1S U29539 ( .I(n24676), .O(n24344) );
  MOAI1S U29540 ( .A1(n24380), .A2(n24680), .B1(n24379), .B2(n24345), .O(
        n24346) );
  INV1S U29541 ( .I(n24407), .O(n24347) );
  NR2 U29542 ( .I1(n24350), .I2(n24347), .O(n24377) );
  MOAI1S U29543 ( .A1(n24472), .A2(n24377), .B1(n24471), .B2(n24348), .O(
        n24349) );
  AOI22S U29544 ( .A1(n24350), .A2(n24484), .B1(n24349), .B2(n24376), .O(
        n24388) );
  INV1S U29545 ( .I(n24351), .O(n24421) );
  NR2 U29546 ( .I1(n24421), .I2(n24418), .O(n24358) );
  INV1S U29547 ( .I(n24353), .O(n24653) );
  ND2S U29548 ( .I1(n24382), .I2(n24654), .O(n24356) );
  ND2S U29549 ( .I1(n24379), .I2(n24354), .O(n24355) );
  ND2S U29550 ( .I1(n24418), .I2(n24421), .O(n24357) );
  OAI12HS U29551 ( .B1(n24358), .B2(n15985), .A1(n24357), .O(n24369) );
  MOAI1 U29552 ( .A1(n24380), .A2(n24646), .B1(n24379), .B2(n24644), .O(n24360) );
  NR2 U29553 ( .I1(n24454), .I2(n15923), .O(n24366) );
  INV1S U29554 ( .I(n24361), .O(n24441) );
  AO12 U29555 ( .B1(n24382), .B2(n24640), .A1(n24362), .O(n24440) );
  NR2 U29556 ( .I1(n24441), .I2(n24440), .O(n24363) );
  NR2 U29557 ( .I1(n24366), .I2(n24363), .O(n24368) );
  ND2S U29558 ( .I1(n24440), .I2(n24441), .O(n24365) );
  ND2S U29559 ( .I1(n15923), .I2(n24454), .O(n24364) );
  OAI12HS U29560 ( .B1(n24366), .B2(n24365), .A1(n24364), .O(n24367) );
  AOI12HS U29561 ( .B1(n24369), .B2(n24368), .A1(n24367), .O(n24374) );
  INV1S U29562 ( .I(n24370), .O(n24496) );
  NR2 U29563 ( .I1(n24496), .I2(n24495), .O(n24373) );
  ND2S U29564 ( .I1(n24495), .I2(n24496), .O(n24372) );
  OAI12HS U29565 ( .B1(n24374), .B2(n24373), .A1(n24372), .O(n24383) );
  INV1S U29566 ( .I(n24375), .O(n24509) );
  ND2S U29567 ( .I1(n24383), .I2(n24509), .O(n24386) );
  INV1S U29568 ( .I(n24376), .O(n24473) );
  AOI12HS U29569 ( .B1(n24472), .B2(n24473), .A1(n24377), .O(n24385) );
  MOAI1S U29570 ( .A1(n24380), .A2(n24696), .B1(n24379), .B2(n24378), .O(
        n24381) );
  OAI12HS U29571 ( .B1(n24383), .B2(n24509), .A1(n24508), .O(n24384) );
  ND3HT U29572 ( .I1(n24389), .I2(n24388), .I3(n24387), .O(n24759) );
  NR2 U29573 ( .I1(n24452), .I2(n15923), .O(n24395) );
  NR2 U29574 ( .I1(n24439), .I2(n24440), .O(n24390) );
  NR2 U29575 ( .I1(n24395), .I2(n24390), .O(n24398) );
  NR2 U29576 ( .I1(n24417), .I2(n24418), .O(n24392) );
  ND2S U29577 ( .I1(n24418), .I2(n24417), .O(n24391) );
  OAI12HS U29578 ( .B1(n24392), .B2(n15985), .A1(n24391), .O(n24397) );
  ND2S U29579 ( .I1(n24440), .I2(n24439), .O(n24394) );
  ND2S U29580 ( .I1(n15923), .I2(n24452), .O(n24393) );
  OAI12HS U29581 ( .B1(n24395), .B2(n24394), .A1(n24393), .O(n24396) );
  AOI12HS U29582 ( .B1(n24398), .B2(n24397), .A1(n24396), .O(n24416) );
  NR2 U29583 ( .I1(n24507), .I2(n24508), .O(n24405) );
  NR2 U29584 ( .I1(n24494), .I2(n24495), .O(n24399) );
  NR2 U29585 ( .I1(n24405), .I2(n24399), .O(n24402) );
  INV1S U29586 ( .I(n24400), .O(n24406) );
  NR2 U29587 ( .I1(n24406), .I2(n24407), .O(n24409) );
  NR2 U29588 ( .I1(n24471), .I2(n24472), .O(n24401) );
  NR2 U29589 ( .I1(n24409), .I2(n24401), .O(n24413) );
  ND2S U29590 ( .I1(n24402), .I2(n24413), .O(n24415) );
  ND2S U29591 ( .I1(n24495), .I2(n24494), .O(n24404) );
  ND2S U29592 ( .I1(n24508), .I2(n24507), .O(n24403) );
  OAI12HS U29593 ( .B1(n24405), .B2(n24404), .A1(n24403), .O(n24412) );
  ND2S U29594 ( .I1(n24472), .I2(n24471), .O(n24410) );
  ND2S U29595 ( .I1(n24407), .I2(n24406), .O(n24408) );
  OAI12HS U29596 ( .B1(n24410), .B2(n24409), .A1(n24408), .O(n24411) );
  AOI12HS U29597 ( .B1(n24413), .B2(n24412), .A1(n24411), .O(n24414) );
  OAI12HS U29598 ( .B1(n24416), .B2(n24415), .A1(n24414), .O(n24419) );
  ND2P U29599 ( .I1(n24759), .I2(n24419), .O(n24770) );
  NR2 U29600 ( .I1(n24417), .I2(n24770), .O(n24424) );
  INV1S U29601 ( .I(n24418), .O(n24422) );
  INV1S U29602 ( .I(n24419), .O(n24420) );
  OAI22S U29603 ( .A1(n24422), .A2(n24758), .B1(n24421), .B2(n24759), .O(
        n24423) );
  ND2S U29604 ( .I1(n24514), .I2(n24425), .O(n24438) );
  ND2S U29605 ( .I1(n24517), .I2(n24426), .O(n24437) );
  INV1S U29606 ( .I(n24610), .O(n24860) );
  INV1S U29607 ( .I(n24763), .O(n24428) );
  ND3S U29608 ( .I1(n24860), .I2(n24428), .I3(n24762), .O(n24433) );
  INV1S U29609 ( .I(n24608), .O(n24858) );
  ND3S U29610 ( .I1(n24858), .I2(n24431), .I3(n24856), .O(n24432) );
  OAI112HS U29611 ( .C1(n24434), .C2(n24861), .A1(n24433), .B1(n24432), .O(
        n24435) );
  ND2S U29612 ( .I1(n24519), .I2(n24435), .O(n24436) );
  ND3 U29613 ( .I1(n24438), .I2(n24437), .I3(n24436), .O(n24869) );
  MAO222 U29614 ( .A1(n24851), .B1(n24853), .C1(n24869), .O(n24466) );
  NR2 U29615 ( .I1(n24439), .I2(n24770), .O(n24444) );
  INV1S U29616 ( .I(n24440), .O(n24442) );
  OAI22S U29617 ( .A1(n24442), .A2(n24758), .B1(n24441), .B2(n24759), .O(
        n24443) );
  ND2S U29618 ( .I1(n24514), .I2(n24445), .O(n24451) );
  ND2S U29619 ( .I1(n24517), .I2(n24446), .O(n24450) );
  INV1S U29620 ( .I(n24447), .O(n24448) );
  ND2S U29621 ( .I1(n24519), .I2(n24448), .O(n24449) );
  OR2 U29622 ( .I1(n24873), .I2(n24825), .O(n24465) );
  NR2 U29623 ( .I1(n24452), .I2(n24770), .O(n24457) );
  INV1S U29624 ( .I(n15923), .O(n24455) );
  OAI22S U29625 ( .A1(n24455), .A2(n24758), .B1(n24454), .B2(n24759), .O(
        n24456) );
  NR2P U29626 ( .I1(n24457), .I2(n24456), .O(n24876) );
  INV1S U29627 ( .I(n24458), .O(n24459) );
  ND2S U29628 ( .I1(n24519), .I2(n24459), .O(n24464) );
  ND2S U29629 ( .I1(n24517), .I2(n24460), .O(n24463) );
  ND2S U29630 ( .I1(n24514), .I2(n24461), .O(n24462) );
  OR2 U29631 ( .I1(n24876), .I2(n24828), .O(n24467) );
  ND3 U29632 ( .I1(n24466), .I2(n24465), .I3(n24467), .O(n24470) );
  ND2S U29633 ( .I1(n24828), .I2(n24876), .O(n24468) );
  ND3 U29634 ( .I1(n24470), .I2(n24469), .I3(n24468), .O(n24525) );
  NR2 U29635 ( .I1(n24471), .I2(n24770), .O(n24476) );
  INV1S U29636 ( .I(n24472), .O(n24474) );
  OAI22S U29637 ( .A1(n24474), .A2(n24758), .B1(n24473), .B2(n24759), .O(
        n24475) );
  ND2S U29638 ( .I1(n24514), .I2(n24477), .O(n24483) );
  INV1S U29639 ( .I(n24478), .O(n24479) );
  ND2S U29640 ( .I1(n24517), .I2(n24479), .O(n24482) );
  ND2S U29641 ( .I1(n24519), .I2(n24480), .O(n24481) );
  NR2 U29642 ( .I1(n24888), .I2(n24887), .O(n24493) );
  ND2S U29643 ( .I1(n24514), .I2(n24486), .O(n24492) );
  INV1S U29644 ( .I(n24487), .O(n24488) );
  ND2S U29645 ( .I1(n24517), .I2(n24488), .O(n24491) );
  ND2S U29646 ( .I1(n24519), .I2(n24489), .O(n24490) );
  NR2 U29647 ( .I1(n24894), .I2(n24817), .O(n24526) );
  NR2 U29648 ( .I1(n24493), .I2(n24526), .O(n24532) );
  NR2 U29649 ( .I1(n24494), .I2(n24770), .O(n24499) );
  INV1S U29650 ( .I(n24495), .O(n24497) );
  OAI22S U29651 ( .A1(n24497), .A2(n24758), .B1(n24496), .B2(n24759), .O(
        n24498) );
  NR2 U29652 ( .I1(n24499), .I2(n24498), .O(n24880) );
  ND2S U29653 ( .I1(n24514), .I2(n24500), .O(n24506) );
  INV1S U29654 ( .I(n24501), .O(n24502) );
  ND2S U29655 ( .I1(n24517), .I2(n24502), .O(n24505) );
  ND2S U29656 ( .I1(n24519), .I2(n24503), .O(n24504) );
  ND3 U29657 ( .I1(n24506), .I2(n24505), .I3(n24504), .O(n24820) );
  NR2 U29658 ( .I1(n24880), .I2(n24820), .O(n24523) );
  NR2 U29659 ( .I1(n24507), .I2(n24770), .O(n24512) );
  INV1S U29660 ( .I(n24508), .O(n24510) );
  OAI22S U29661 ( .A1(n24510), .A2(n24758), .B1(n24509), .B2(n24759), .O(
        n24511) );
  NR2 U29662 ( .I1(n24512), .I2(n24511), .O(n24884) );
  ND2S U29663 ( .I1(n24514), .I2(n24513), .O(n24522) );
  INV1S U29664 ( .I(n24515), .O(n24516) );
  ND2S U29665 ( .I1(n24517), .I2(n24516), .O(n24521) );
  ND2S U29666 ( .I1(n24519), .I2(n24518), .O(n24520) );
  NR2 U29667 ( .I1(n24884), .I2(n24819), .O(n24531) );
  NR2 U29668 ( .I1(n24523), .I2(n24531), .O(n24524) );
  ND3 U29669 ( .I1(n24525), .I2(n24532), .I3(n24524), .O(n24536) );
  INV1S U29670 ( .I(n24526), .O(n24529) );
  INV1S U29671 ( .I(n24894), .O(n24527) );
  INV1S U29672 ( .I(n24817), .O(n24891) );
  NR2 U29673 ( .I1(n24527), .I2(n24891), .O(n24528) );
  AOI13HS U29674 ( .B1(n24529), .B2(n24888), .B3(n24887), .A1(n24528), .O(
        n24535) );
  ND2S U29675 ( .I1(n24820), .I2(n24880), .O(n24530) );
  MOAI1 U29676 ( .A1(n24531), .A2(n24530), .B1(n24819), .B2(n24884), .O(n24533) );
  ND2S U29677 ( .I1(n24533), .I2(n24532), .O(n24534) );
  ND3P U29678 ( .I1(n24536), .I2(n24535), .I3(n24534), .O(n24849) );
  INV1S U29679 ( .I(n24604), .O(n24620) );
  ND2S U29680 ( .I1(n24614), .I2(mem_data_out_reg_shift_1[19]), .O(n24539) );
  ND2S U29681 ( .I1(n24616), .I2(n24537), .O(n24538) );
  ND2S U29682 ( .I1(n24608), .I2(n24541), .O(n24544) );
  ND2S U29683 ( .I1(n24610), .I2(n24542), .O(n24543) );
  OAI112HS U29684 ( .C1(n24862), .C2(n24545), .A1(n24544), .B1(n24543), .O(
        n24743) );
  NR2 U29685 ( .I1(n24743), .I2(n24747), .O(n24574) );
  ND2S U29686 ( .I1(n24608), .I2(n24546), .O(n24549) );
  ND2S U29687 ( .I1(n24610), .I2(n24547), .O(n24548) );
  OAI112HS U29688 ( .C1(n24862), .C2(n24550), .A1(n24549), .B1(n24548), .O(
        n24748) );
  BUF1S U29689 ( .I(n24614), .O(n24583) );
  ND2S U29690 ( .I1(n24583), .I2(mem_data_out_reg_shift_1[18]), .O(n24553) );
  ND2S U29691 ( .I1(n24616), .I2(n24551), .O(n24552) );
  NR2 U29692 ( .I1(n24748), .I2(n24752), .O(n24555) );
  NR2 U29693 ( .I1(n24574), .I2(n24555), .O(n24577) );
  ND2S U29694 ( .I1(n24610), .I2(n24556), .O(n24559) );
  ND2S U29695 ( .I1(n24608), .I2(n24557), .O(n24558) );
  OAI112HS U29696 ( .C1(n24862), .C2(n24560), .A1(n24559), .B1(n24558), .O(
        n24757) );
  INV1S U29697 ( .I(n24561), .O(n24565) );
  ND2S U29698 ( .I1(n24616), .I2(n24562), .O(n24564) );
  ND2S U29699 ( .I1(n24583), .I2(mem_data_out_reg_shift_1[16]), .O(n24563) );
  NR2 U29700 ( .I1(n24757), .I2(n24867), .O(n24571) );
  ND2S U29701 ( .I1(n24614), .I2(mem_data_out_reg_shift_1[17]), .O(n24568) );
  ND2S U29702 ( .I1(n24616), .I2(n24566), .O(n24567) );
  OAI112HS U29703 ( .C1(n24620), .C2(n24569), .A1(n24568), .B1(n24567), .O(
        n24754) );
  ND2S U29704 ( .I1(n24867), .I2(n24757), .O(n24570) );
  OAI12HS U29705 ( .B1(n24571), .B2(n24754), .A1(n24570), .O(n24576) );
  ND2S U29706 ( .I1(n24752), .I2(n24748), .O(n24573) );
  ND2S U29707 ( .I1(n24747), .I2(n24743), .O(n24572) );
  OAI12HS U29708 ( .B1(n24574), .B2(n24573), .A1(n24572), .O(n24575) );
  AOI12HS U29709 ( .B1(n24577), .B2(n24576), .A1(n24575), .O(n24635) );
  ND2S U29710 ( .I1(n24608), .I2(n24578), .O(n24581) );
  ND2S U29711 ( .I1(n24610), .I2(n24579), .O(n24580) );
  OAI112HS U29712 ( .C1(n24862), .C2(n24582), .A1(n24581), .B1(n24580), .O(
        n24786) );
  ND2S U29713 ( .I1(n24583), .I2(mem_data_out_reg_shift_1[20]), .O(n24586) );
  ND2S U29714 ( .I1(n24616), .I2(n24584), .O(n24585) );
  NR2 U29715 ( .I1(n24786), .I2(n24790), .O(n24597) );
  ND2S U29716 ( .I1(n24608), .I2(n24588), .O(n24591) );
  ND2S U29717 ( .I1(n24610), .I2(n24589), .O(n24590) );
  OAI112HS U29718 ( .C1(n24862), .C2(n24592), .A1(n24591), .B1(n24590), .O(
        n24781) );
  ND2S U29719 ( .I1(n24614), .I2(mem_data_out_reg_shift_1[21]), .O(n24595) );
  ND2S U29720 ( .I1(n24616), .I2(n24593), .O(n24594) );
  NR2 U29721 ( .I1(n24781), .I2(n24785), .O(n24625) );
  NR2 U29722 ( .I1(n24597), .I2(n24625), .O(n24622) );
  ND3S U29723 ( .I1(n24600), .I2(n24599), .I3(n24598), .O(n24792) );
  INV1S U29724 ( .I(n24792), .O(n24626) );
  ND2S U29725 ( .I1(n24601), .I2(mem_data_out_reg_shift_1[23]), .O(n24603) );
  ND2S U29726 ( .I1(n24603), .I2(n24602), .O(n24606) );
  MXL2HS U29727 ( .A(n24606), .B(n24605), .S(n24604), .OB(n24793) );
  NR2 U29728 ( .I1(n24626), .I2(n24793), .O(n24628) );
  ND2S U29729 ( .I1(n24608), .I2(n24607), .O(n24612) );
  ND2S U29730 ( .I1(n24610), .I2(n24609), .O(n24611) );
  OAI112HS U29731 ( .C1(n24862), .C2(n24613), .A1(n24612), .B1(n24611), .O(
        n24796) );
  ND2S U29732 ( .I1(n24614), .I2(mem_data_out_reg_shift_1[22]), .O(n24618) );
  ND2S U29733 ( .I1(n24616), .I2(n24615), .O(n24617) );
  NR2 U29734 ( .I1(n24796), .I2(n24801), .O(n24621) );
  NR2 U29735 ( .I1(n24628), .I2(n24621), .O(n24631) );
  ND2S U29736 ( .I1(n24622), .I2(n24631), .O(n24634) );
  ND2S U29737 ( .I1(n24790), .I2(n24786), .O(n24624) );
  ND2S U29738 ( .I1(n24785), .I2(n24781), .O(n24623) );
  OAI12HS U29739 ( .B1(n24625), .B2(n24624), .A1(n24623), .O(n24632) );
  ND2S U29740 ( .I1(n24801), .I2(n24796), .O(n24629) );
  ND2S U29741 ( .I1(n24793), .I2(n24626), .O(n24627) );
  OAI12HS U29742 ( .B1(n24629), .B2(n24628), .A1(n24627), .O(n24630) );
  AOI12HS U29743 ( .B1(n24632), .B2(n24631), .A1(n24630), .O(n24633) );
  OAI12HS U29744 ( .B1(n24635), .B2(n24634), .A1(n24633), .O(n24716) );
  INV1S U29745 ( .I(n24636), .O(n24637) );
  ND2S U29746 ( .I1(n24698), .I2(n24640), .O(n24641) );
  NR2 U29747 ( .I1(n24752), .I2(n24749), .O(n24651) );
  INV1S U29748 ( .I(n24644), .O(n24645) );
  OR2 U29749 ( .I1(n24645), .I2(n24693), .O(n24650) );
  OR2 U29750 ( .I1(n24646), .I2(n24695), .O(n24649) );
  ND2S U29751 ( .I1(n24698), .I2(n24647), .O(n24648) );
  ND3P U29752 ( .I1(n24650), .I2(n24649), .I3(n24648), .O(n24744) );
  NR2 U29753 ( .I1(n24747), .I2(n24744), .O(n24670) );
  NR2 U29754 ( .I1(n24651), .I2(n24670), .O(n24673) );
  ND2S U29755 ( .I1(n24698), .I2(n24654), .O(n24655) );
  ND3S U29756 ( .I1(n24657), .I2(n24656), .I3(n24655), .O(n24718) );
  NR2 U29757 ( .I1(n24665), .I2(n24718), .O(n24667) );
  INV1S U29758 ( .I(n24658), .O(n24659) );
  ND2S U29759 ( .I1(n24698), .I2(n24661), .O(n24662) );
  ND2S U29760 ( .I1(n24718), .I2(n24665), .O(n24666) );
  OAI12HS U29761 ( .B1(n24667), .B2(n15984), .A1(n24666), .O(n24672) );
  ND2S U29762 ( .I1(n24749), .I2(n24752), .O(n24669) );
  ND2S U29763 ( .I1(n24744), .I2(n24747), .O(n24668) );
  OAI12HS U29764 ( .B1(n24670), .B2(n24669), .A1(n24668), .O(n24671) );
  AOI12HS U29765 ( .B1(n24673), .B2(n24672), .A1(n24671), .O(n24715) );
  INV1S U29766 ( .I(n24674), .O(n24675) );
  ND2S U29767 ( .I1(n24676), .I2(n24675), .O(n24678) );
  MXL2HS U29768 ( .A(n24678), .B(n24677), .S(n24698), .OB(n24794) );
  NR2 U29769 ( .I1(n24793), .I2(n24794), .O(n24708) );
  ND2S U29770 ( .I1(n24698), .I2(n24681), .O(n24682) );
  ND3 U29771 ( .I1(n24684), .I2(n24683), .I3(n24682), .O(n24797) );
  NR2 U29772 ( .I1(n24801), .I2(n24797), .O(n24685) );
  NR2 U29773 ( .I1(n24708), .I2(n24685), .O(n24712) );
  INV1S U29774 ( .I(n24686), .O(n24687) );
  ND2S U29775 ( .I1(n24698), .I2(n24689), .O(n24690) );
  ND3S U29776 ( .I1(n24692), .I2(n24691), .I3(n24690), .O(n24787) );
  NR2 U29777 ( .I1(n24790), .I2(n24787), .O(n24702) );
  ND2S U29778 ( .I1(n24698), .I2(n24697), .O(n24699) );
  ND3S U29779 ( .I1(n24701), .I2(n24700), .I3(n24699), .O(n24782) );
  NR2 U29780 ( .I1(n24785), .I2(n24782), .O(n24706) );
  NR2 U29781 ( .I1(n24702), .I2(n24706), .O(n24703) );
  ND2S U29782 ( .I1(n24712), .I2(n24703), .O(n24714) );
  ND2S U29783 ( .I1(n24787), .I2(n24790), .O(n24705) );
  ND2S U29784 ( .I1(n24782), .I2(n24785), .O(n24704) );
  OAI12HS U29785 ( .B1(n24706), .B2(n24705), .A1(n24704), .O(n24711) );
  ND2S U29786 ( .I1(n24797), .I2(n24801), .O(n24709) );
  OAI12HS U29787 ( .B1(n24709), .B2(n24708), .A1(n24707), .O(n24710) );
  AOI12HS U29788 ( .B1(n24712), .B2(n24711), .A1(n24710), .O(n24713) );
  OAI12HS U29789 ( .B1(n24715), .B2(n24714), .A1(n24713), .O(n24739) );
  NR2P U29790 ( .I1(n24716), .I2(n24739), .O(n24755) );
  INV1S U29791 ( .I(n24744), .O(n24722) );
  NR2 U29792 ( .I1(n24743), .I2(n24722), .O(n24725) );
  INV1S U29793 ( .I(n24749), .O(n24721) );
  NR2 U29794 ( .I1(n24748), .I2(n24721), .O(n24717) );
  NR2 U29795 ( .I1(n24725), .I2(n24717), .O(n24728) );
  NR2 U29796 ( .I1(n24757), .I2(n15984), .O(n24720) );
  INV1S U29797 ( .I(n24718), .O(n24865) );
  ND2S U29798 ( .I1(n15984), .I2(n24757), .O(n24719) );
  OAI12HS U29799 ( .B1(n24720), .B2(n24718), .A1(n24719), .O(n24727) );
  ND2S U29800 ( .I1(n24721), .I2(n24748), .O(n24724) );
  ND2S U29801 ( .I1(n24722), .I2(n24743), .O(n24723) );
  OAI12HS U29802 ( .B1(n24725), .B2(n24724), .A1(n24723), .O(n24726) );
  AOI12HS U29803 ( .B1(n24728), .B2(n24727), .A1(n24726), .O(n24732) );
  INV1S U29804 ( .I(n24787), .O(n24729) );
  NR2 U29805 ( .I1(n24786), .I2(n24729), .O(n24731) );
  ND2S U29806 ( .I1(n24729), .I2(n24786), .O(n24730) );
  INV1S U29807 ( .I(n24782), .O(n24733) );
  AOI12HS U29808 ( .B1(n24734), .B2(n24781), .A1(n24733), .O(n24737) );
  NR2 U29809 ( .I1(n24781), .I2(n24734), .O(n24736) );
  INV1S U29810 ( .I(n24797), .O(n24735) );
  MOAI1 U29811 ( .A1(n24737), .A2(n24736), .B1(n24735), .B2(n24796), .O(n24742) );
  INV1S U29812 ( .I(n24796), .O(n24738) );
  AOI22S U29813 ( .A1(n24794), .A2(n24792), .B1(n24797), .B2(n24738), .O(
        n24741) );
  OAI12HS U29814 ( .B1(n24794), .B2(n24792), .A1(n24739), .O(n24740) );
  AOI12H U29815 ( .B1(n24742), .B2(n24741), .A1(n24740), .O(n24798) );
  ND2S U29816 ( .I1(n24855), .I2(n24743), .O(n24746) );
  ND2S U29817 ( .I1(n24798), .I2(n24744), .O(n24745) );
  OAI112HS U29818 ( .C1(n24747), .C2(n24868), .A1(n24746), .B1(n24745), .O(
        n24827) );
  NR2 U29819 ( .I1(n24876), .I2(n24827), .O(n24777) );
  ND2S U29820 ( .I1(n24855), .I2(n24748), .O(n24751) );
  ND2S U29821 ( .I1(n24798), .I2(n24749), .O(n24750) );
  OAI112HS U29822 ( .C1(n24752), .C2(n24868), .A1(n24751), .B1(n24750), .O(
        n24824) );
  NR2 U29823 ( .I1(n24873), .I2(n24824), .O(n24753) );
  NR2 U29824 ( .I1(n24777), .I2(n24753), .O(n24780) );
  INV1S U29825 ( .I(n24798), .O(n24866) );
  MOAI1S U29826 ( .A1(n24866), .A2(n15984), .B1(n24755), .B2(n24754), .O(
        n24756) );
  AOI12HS U29827 ( .B1(n24855), .B2(n24757), .A1(n24756), .O(n24854) );
  NR2 U29828 ( .I1(n15985), .I2(n24758), .O(n24772) );
  INV1S U29829 ( .I(n24759), .O(n24768) );
  ND2S U29830 ( .I1(n24761), .I2(n24760), .O(n24766) );
  AOI22S U29831 ( .A1(n24764), .A2(n24856), .B1(n24763), .B2(n24762), .O(
        n24765) );
  ND2S U29832 ( .I1(n24766), .I2(n24765), .O(n24767) );
  MOAI1S U29833 ( .A1(n24770), .A2(n24769), .B1(n24768), .B2(n24767), .O(
        n24771) );
  NR2 U29834 ( .I1(n24870), .I2(n24853), .O(n24774) );
  ND2S U29835 ( .I1(n24853), .I2(n24870), .O(n24773) );
  OAI12HS U29836 ( .B1(n24854), .B2(n24774), .A1(n24773), .O(n24779) );
  ND2S U29837 ( .I1(n24824), .I2(n24873), .O(n24776) );
  ND2S U29838 ( .I1(n24827), .I2(n24876), .O(n24775) );
  OAI12HS U29839 ( .B1(n24777), .B2(n24776), .A1(n24775), .O(n24778) );
  AOI12HS U29840 ( .B1(n24780), .B2(n24779), .A1(n24778), .O(n24815) );
  ND2S U29841 ( .I1(n24855), .I2(n24781), .O(n24784) );
  ND2S U29842 ( .I1(n24798), .I2(n24782), .O(n24783) );
  NR2 U29843 ( .I1(n24884), .I2(n24883), .O(n24806) );
  ND2S U29844 ( .I1(n24855), .I2(n24786), .O(n24789) );
  ND2S U29845 ( .I1(n24798), .I2(n24787), .O(n24788) );
  OAI112HS U29846 ( .C1(n24790), .C2(n24868), .A1(n24789), .B1(n24788), .O(
        n24879) );
  NR2 U29847 ( .I1(n24880), .I2(n24879), .O(n24791) );
  NR2 U29848 ( .I1(n24806), .I2(n24791), .O(n24803) );
  ND2S U29849 ( .I1(n24793), .I2(n24792), .O(n24795) );
  NR2 U29850 ( .I1(n24894), .I2(n24835), .O(n24808) );
  ND2S U29851 ( .I1(n24798), .I2(n24797), .O(n24799) );
  NR2 U29852 ( .I1(n24888), .I2(n24816), .O(n24802) );
  NR2 U29853 ( .I1(n24808), .I2(n24802), .O(n24811) );
  ND2S U29854 ( .I1(n24803), .I2(n24811), .O(n24814) );
  ND2S U29855 ( .I1(n24879), .I2(n24880), .O(n24805) );
  ND2S U29856 ( .I1(n24883), .I2(n24884), .O(n24804) );
  OAI12HS U29857 ( .B1(n24806), .B2(n24805), .A1(n24804), .O(n24812) );
  ND2S U29858 ( .I1(n24816), .I2(n24888), .O(n24809) );
  OAI12HS U29859 ( .B1(n24809), .B2(n24808), .A1(n24807), .O(n24810) );
  AOI12HS U29860 ( .B1(n24812), .B2(n24811), .A1(n24810), .O(n24813) );
  OAI12HS U29861 ( .B1(n24815), .B2(n24814), .A1(n24813), .O(n24844) );
  INV3CK U29862 ( .I(n24816), .O(n24890) );
  NR2 U29863 ( .I1(n24890), .I2(n24887), .O(n24818) );
  INV1S U29864 ( .I(n24835), .O(n24895) );
  NR2 U29865 ( .I1(n24895), .I2(n24817), .O(n24836) );
  NR2 U29866 ( .I1(n24818), .I2(n24836), .O(n24841) );
  ND2S U29867 ( .I1(n24885), .I2(n24883), .O(n24830) );
  INV1S U29868 ( .I(n24820), .O(n24881) );
  NR2 U29869 ( .I1(n24879), .I2(n24881), .O(n24821) );
  MOAI1 U29870 ( .A1(n24885), .A2(n24883), .B1(n24830), .B2(n24821), .O(n24840) );
  INV1S U29871 ( .I(n24825), .O(n24874) );
  ND2S U29872 ( .I1(n24874), .I2(n24824), .O(n24823) );
  INV1S U29873 ( .I(n24828), .O(n24877) );
  ND2S U29874 ( .I1(n24877), .I2(n24827), .O(n24826) );
  MAO222 U29875 ( .A1(n24869), .B1(n24854), .C1(n24851), .O(n24822) );
  ND3S U29876 ( .I1(n24823), .I2(n24826), .I3(n24822), .O(n24834) );
  INV1S U29877 ( .I(n24824), .O(n24875) );
  ND3S U29878 ( .I1(n24826), .I2(n24875), .I3(n24825), .O(n24833) );
  INV1S U29879 ( .I(n24827), .O(n24878) );
  ND2S U29880 ( .I1(n24828), .I2(n24878), .O(n24832) );
  ND2S U29881 ( .I1(n24881), .I2(n24879), .O(n24829) );
  ND3 U29882 ( .I1(n24841), .I2(n24830), .I3(n24829), .O(n24831) );
  AOI13HS U29883 ( .B1(n24834), .B2(n24833), .B3(n24832), .A1(n24831), .O(
        n24839) );
  ND2S U29884 ( .I1(n24887), .I2(n24890), .O(n24837) );
  OAI22S U29885 ( .A1(n24837), .A2(n24836), .B1(n24891), .B2(n24835), .O(
        n24838) );
  AO112P U29886 ( .C1(n24841), .C2(n24840), .A1(n24839), .B1(n24838), .O(
        n24848) );
  MUX2 U29887 ( .A(n24850), .B(n24844), .S(n24848), .O(n24842) );
  ND2 U29888 ( .I1(n24850), .I2(n24844), .O(n24843) );
  INV3CK U29889 ( .I(n24843), .O(n24847) );
  INV1S U29890 ( .I(n24844), .O(n24845) );
  AN2 U29891 ( .I1(n24849), .I2(n24845), .O(n24846) );
  NR2F U29892 ( .I1(n24847), .I2(n24846), .O(n24893) );
  MUX2T U29893 ( .A(n24850), .B(n24849), .S(n24848), .O(n24892) );
  INV1S U29894 ( .I(n24851), .O(n24852) );
  OAI222S U29895 ( .A1(n24896), .A2(n24854), .B1(n24853), .B2(n24893), .C1(
        n24892), .C2(n24852), .O(n15858) );
  INV1S U29896 ( .I(n24855), .O(n24864) );
  INV1S U29897 ( .I(n24856), .O(n24857) );
  OA222S U29898 ( .A1(n24862), .A2(n24861), .B1(n24860), .B2(n24859), .C1(
        n24858), .C2(n24857), .O(n24863) );
  INV1S U29899 ( .I(n24869), .O(n24871) );
  OAI222S U29900 ( .A1(n24896), .A2(n24872), .B1(n24871), .B2(n24892), .C1(
        n24870), .C2(n24893), .O(n15857) );
  OAI222S U29901 ( .A1(n24896), .A2(n24875), .B1(n24874), .B2(n24892), .C1(
        n24893), .C2(n24873), .O(n15859) );
  OAI222S U29902 ( .A1(n24896), .A2(n24878), .B1(n24877), .B2(n24892), .C1(
        n24893), .C2(n24876), .O(n15860) );
  INV1S U29903 ( .I(n24879), .O(n24882) );
  OAI222S U29904 ( .A1(n24896), .A2(n24882), .B1(n24881), .B2(n24892), .C1(
        n24893), .C2(n24880), .O(n15861) );
  INV1S U29905 ( .I(n24883), .O(n24886) );
  OAI222S U29906 ( .A1(n24896), .A2(n24886), .B1(n24885), .B2(n24892), .C1(
        n24893), .C2(n24884), .O(n15862) );
  INV1S U29907 ( .I(n24887), .O(n24889) );
  OAI222S U29908 ( .A1(n24896), .A2(n24890), .B1(n24889), .B2(n24892), .C1(
        n24893), .C2(n24888), .O(n15863) );
  OAI222S U29909 ( .A1(n24896), .A2(n24895), .B1(n24894), .B2(n24893), .C1(
        n24892), .C2(n24891), .O(n15864) );
  OAI12HS U29910 ( .B1(n24934), .B2(n24898), .A1(n24897), .O(n15755) );
  INV1S U29911 ( .I(image_size_reg_master[1]), .O(n30394) );
  OAI22S U29912 ( .A1(n24900), .A2(n24899), .B1(n30394), .B2(n30391), .O(
        n15757) );
  MOAI1S U29913 ( .A1(n30412), .A2(n24902), .B1(n30411), .B2(n24901), .O(
        n15754) );
  MOAI1S U29914 ( .A1(n30412), .A2(n24903), .B1(n30411), .B2(
        image_size_reg_set[1]), .O(n15753) );
  XNR2HS U29915 ( .I1(cnt_dyn_base[1]), .I2(medfilt_cnt[1]), .O(n24904) );
  ND3S U29916 ( .I1(n24906), .I2(n24905), .I3(n24904), .O(n24908) );
  OR2S U29917 ( .I1(n24908), .I2(n24907), .O(n30239) );
  MOAI1S U29918 ( .A1(n24910), .A2(cs[1]), .B1(n24909), .B2(medfilt_state[3]), 
        .O(n30238) );
  NR2 U29919 ( .I1(n30239), .I2(n30238), .O(n30425) );
  ND2S U29920 ( .I1(n30425), .I2(medfilt_cnt2[0]), .O(n24912) );
  ND2S U29921 ( .I1(n24912), .I2(medfilt_cnt2[1]), .O(n24911) );
  OAI22S U29922 ( .A1(medfilt_cnt2[1]), .A2(n24912), .B1(n24911), .B2(n30238), 
        .O(n15735) );
  INV1S U29923 ( .I(medfilt_cnt2[1]), .O(n24913) );
  NR2 U29924 ( .I1(n24913), .I2(n24912), .O(n24915) );
  ND2S U29925 ( .I1(medfilt_cnt2[2]), .I2(n24915), .O(n24916) );
  ND2S U29926 ( .I1(n24916), .I2(medfilt_cnt2[3]), .O(n24914) );
  OAI22S U29927 ( .A1(n24914), .A2(n30238), .B1(medfilt_cnt2[3]), .B2(n24916), 
        .O(n15733) );
  ND2S U29928 ( .I1(medfilt_cnt2[2]), .I2(n24916), .O(n24917) );
  MOAI1S U29929 ( .A1(n30238), .A2(n24917), .B1(n24916), .B2(n24915), .O(
        n15734) );
  INV1S U29930 ( .I(n24918), .O(n24920) );
  ND2S U29931 ( .I1(n24920), .I2(n24919), .O(n24926) );
  INV1S U29932 ( .I(n30241), .O(n24921) );
  OAI112HS U29933 ( .C1(n24923), .C2(n24922), .A1(n24932), .B1(n24921), .O(
        n24924) );
  MOAI1S U29934 ( .A1(n30360), .A2(n24926), .B1(n24925), .B2(n24924), .O(N7421) );
  INV1S U29935 ( .I(n24927), .O(n24933) );
  ND2S U29936 ( .I1(n24929), .I2(n24928), .O(n24931) );
  AOI13HS U29937 ( .B1(n24933), .B2(n24932), .B3(n24931), .A1(n24930), .O(
        N7422) );
  NR2 U29938 ( .I1(n24934), .I2(n30371), .O(n24937) );
  INV1S U29939 ( .I(n30298), .O(n30222) );
  ND2S U29940 ( .I1(n30452), .I2(n30222), .O(n24935) );
  MOAI1S U29941 ( .A1(n30255), .A2(n24936), .B1(n24937), .B2(n24935), .O(
        n15805) );
  INV1S U29942 ( .I(n24937), .O(n30254) );
  NR2 U29943 ( .I1(cnt_dyn[0]), .I2(n30254), .O(cnt_dyn_n[0]) );
  INV1S U29944 ( .I(n25040), .O(n24953) );
  ND2S U29945 ( .I1(n24953), .I2(cnt_cro_3[0]), .O(n24938) );
  OAI22S U29946 ( .A1(n24939), .A2(n24944), .B1(n30360), .B2(n24938), .O(
        n15764) );
  NR2 U29947 ( .I1(n24940), .I2(n25040), .O(n24941) );
  MOAI1S U29948 ( .A1(n24944), .A2(n24943), .B1(n24942), .B2(n24941), .O(
        n15763) );
  INV1S U29949 ( .I(n24949), .O(n24947) );
  INV1S U29950 ( .I(n24950), .O(n24946) );
  OAI22S U29951 ( .A1(n24951), .A2(n24950), .B1(n24949), .B2(n24948), .O(
        n15762) );
  INV1S U29952 ( .I(n24952), .O(n24957) );
  AOI13HS U29953 ( .B1(n24957), .B2(cnt_cro_x[1]), .B3(cnt_cro_x[0]), .A1(
        n25035), .O(n24959) );
  NR3 U29954 ( .I1(cnt_cro_x[2]), .I2(n30375), .I3(n24962), .O(n24960) );
  INV1S U29955 ( .I(cnt_cro_x[0]), .O(n24956) );
  NR2 U29956 ( .I1(cnt_cro_x[0]), .I2(n24953), .O(n24954) );
  MOAI1S U29957 ( .A1(n24957), .A2(n24956), .B1(n24955), .B2(n24954), .O(
        n15752) );
  INV1S U29958 ( .I(n24962), .O(n24958) );
  NR2 U29959 ( .I1(n24960), .I2(n24959), .O(n24963) );
  ND3S U29960 ( .I1(n30374), .I2(cnt_cro_x[2]), .I3(cnt_cro_x[1]), .O(n24961)
         );
  OAI22S U29961 ( .A1(n30374), .A2(n24963), .B1(n24962), .B2(n24961), .O(
        n15749) );
  ND2S U29962 ( .I1(n16006), .I2(action_done), .O(n24964) );
  NR2 U29963 ( .I1(n30409), .I2(n24964), .O(n24965) );
  XNR2HS U29964 ( .I1(action_5_flag), .I2(n24965), .O(n24966) );
  NR2 U29965 ( .I1(n24967), .I2(n24966), .O(n13612) );
  MOAI1S U29966 ( .A1(n25357), .A2(n25066), .B1(n25355), .B2(n25065), .O(
        n24968) );
  NR2 U29967 ( .I1(n15889), .I2(n24968), .O(n25458) );
  INV1S U29968 ( .I(n25458), .O(n25460) );
  MUX2S U29969 ( .A(n27447), .B(n25458), .S(gray_img[1879]), .O(n24969) );
  MOAI1S U29970 ( .A1(n25062), .A2(n25357), .B1(n25061), .B2(n25355), .O(
        n24970) );
  NR2 U29971 ( .I1(n15889), .I2(n24970), .O(n25759) );
  INV1S U29972 ( .I(n25759), .O(n25761) );
  MOAI1S U29973 ( .A1(n25352), .A2(n25066), .B1(n25351), .B2(n25065), .O(
        n24974) );
  NR2 U29974 ( .I1(n27447), .I2(n24974), .O(n25475) );
  ND2S U29975 ( .I1(n25475), .I2(gray_img[1887]), .O(n24977) );
  OAI112HS U29976 ( .C1(n25291), .C2(n25475), .A1(n24977), .B1(n24976), .O(
        n15488) );
  MOAI1S U29977 ( .A1(n25062), .A2(n25352), .B1(n25061), .B2(n25351), .O(
        n24978) );
  NR2 U29978 ( .I1(n15889), .I2(n24978), .O(n25471) );
  INV1S U29979 ( .I(n25471), .O(n25473) );
  INV1S U29980 ( .I(n24981), .O(n24983) );
  ND2S U29981 ( .I1(n24983), .I2(n24982), .O(n24984) );
  AOI22S U29982 ( .A1(n16006), .A2(n24985), .B1(n25315), .B2(n24984), .O(
        n24986) );
  ND2S U29983 ( .I1(n25291), .I2(n24986), .O(n24987) );
  MUX2S U29984 ( .A(gray_img[943]), .B(n24987), .S(n25612), .O(n13817) );
  MOAI1S U29985 ( .A1(n25357), .A2(n25054), .B1(n25355), .B2(n25053), .O(
        n24988) );
  NR2 U29986 ( .I1(n15889), .I2(n24988), .O(n25492) );
  INV1S U29987 ( .I(n25492), .O(n25494) );
  MOAI1S U29988 ( .A1(n25357), .A2(n25058), .B1(n25355), .B2(n25057), .O(
        n24990) );
  NR2 U29989 ( .I1(n15889), .I2(n24990), .O(n25496) );
  INV1S U29990 ( .I(n25496), .O(n25498) );
  MOAI1S U29991 ( .A1(n25352), .A2(n25054), .B1(n25351), .B2(n25053), .O(
        n24992) );
  NR2 U29992 ( .I1(n27447), .I2(n24992), .O(n25574) );
  INV1S U29993 ( .I(n25574), .O(n25576) );
  MOAI1S U29994 ( .A1(n25352), .A2(n25058), .B1(n25351), .B2(n25057), .O(
        n24994) );
  NR2 U29995 ( .I1(n27447), .I2(n24994), .O(n25508) );
  INV1S U29996 ( .I(n25508), .O(n25510) );
  MOAI1S U29997 ( .A1(n25062), .A2(n25366), .B1(n25061), .B2(n25365), .O(
        n25000) );
  NR2 U29998 ( .I1(n27447), .I2(n25000), .O(n28801) );
  INV1S U29999 ( .I(n28801), .O(n28803) );
  MOAI1S U30000 ( .A1(n25366), .A2(n25066), .B1(n25365), .B2(n25065), .O(
        n25003) );
  NR2 U30001 ( .I1(n15889), .I2(n25003), .O(n25629) );
  ND2S U30002 ( .I1(n25629), .I2(gray_img[1871]), .O(n25006) );
  OAI112HS U30003 ( .C1(n25291), .C2(n25629), .A1(n25006), .B1(n25005), .O(
        n15490) );
  INV1S U30004 ( .I(n25007), .O(n25009) );
  ND2S U30005 ( .I1(n25009), .I2(n25008), .O(n25010) );
  AOI22S U30006 ( .A1(n16006), .A2(n25011), .B1(n25315), .B2(n25010), .O(
        n25012) );
  ND2S U30007 ( .I1(n25291), .I2(n25012), .O(n25013) );
  MUX2S U30008 ( .A(gray_img[935]), .B(n25013), .S(n25751), .O(n13820) );
  MOAI1S U30009 ( .A1(n25366), .A2(n25054), .B1(n25365), .B2(n25053), .O(
        n25014) );
  NR2 U30010 ( .I1(n15889), .I2(n25014), .O(n25651) );
  ND2S U30011 ( .I1(n25651), .I2(gray_img[1615]), .O(n25016) );
  ND2S U30012 ( .I1(n27447), .I2(n25666), .O(n25015) );
  OAI112HS U30013 ( .C1(n25291), .C2(n25651), .A1(n25016), .B1(n25015), .O(
        n15522) );
  MOAI1S U30014 ( .A1(n25366), .A2(n25058), .B1(n25365), .B2(n25057), .O(
        n25017) );
  NR2 U30015 ( .I1(n27447), .I2(n25017), .O(n25647) );
  ND2S U30016 ( .I1(n25647), .I2(gray_img[1743]), .O(n25019) );
  INV1S U30017 ( .I(gray_img[1743]), .O(n25020) );
  ND2S U30018 ( .I1(n27447), .I2(n25020), .O(n25018) );
  OAI112HS U30019 ( .C1(n25291), .C2(n25647), .A1(n25019), .B1(n25018), .O(
        n15506) );
  ND2S U30020 ( .I1(n25020), .I2(n25666), .O(n25687) );
  INV1S U30021 ( .I(n25687), .O(n25021) );
  NR2 U30022 ( .I1(gray_img[1607]), .I2(gray_img[1735]), .O(n25686) );
  ND2S U30023 ( .I1(n25021), .I2(n25686), .O(n25022) );
  AOI22S U30024 ( .A1(n16006), .A2(n25023), .B1(n25315), .B2(n25022), .O(
        n25024) );
  ND2S U30025 ( .I1(n25291), .I2(n25024), .O(n25026) );
  AOI22S U30026 ( .A1(n25103), .A2(n25194), .B1(n25356), .B2(n25193), .O(
        n25025) );
  MUX2S U30027 ( .A(gray_img[807]), .B(n25026), .S(n25744), .O(n13878) );
  INV1S U30028 ( .I(n25027), .O(n25029) );
  ND2S U30029 ( .I1(n25029), .I2(n25028), .O(n25030) );
  AOI22S U30030 ( .A1(n16006), .A2(n28746), .B1(n25315), .B2(n25030), .O(
        n25031) );
  ND2S U30031 ( .I1(n25291), .I2(n25031), .O(n25032) );
  MUX2S U30032 ( .A(gray_img[407]), .B(n25032), .S(n28807), .O(n13616) );
  NR2 U30033 ( .I1(n25037), .I2(n25038), .O(n25042) );
  INV1S U30034 ( .I(n25041), .O(n25033) );
  NR2 U30035 ( .I1(n25042), .I2(n25033), .O(n25036) );
  NR2 U30036 ( .I1(n25036), .I2(n25047), .O(n25044) );
  NR2 U30037 ( .I1(n25044), .I2(n25039), .O(n15746) );
  ND2S U30038 ( .I1(n25042), .I2(n25045), .O(n25043) );
  OAI22S U30039 ( .A1(n25045), .A2(n25044), .B1(n25046), .B2(n25043), .O(
        n15745) );
  INV1S U30040 ( .I(n25046), .O(n25048) );
  MOAI1S U30041 ( .A1(n25341), .A2(n25054), .B1(n25339), .B2(n25053), .O(
        n25055) );
  NR2 U30042 ( .I1(n15889), .I2(n25055), .O(n25897) );
  INV1S U30043 ( .I(n25897), .O(n25899) );
  MOAI1S U30044 ( .A1(n25341), .A2(n25058), .B1(n25339), .B2(n25057), .O(
        n25059) );
  NR2 U30045 ( .I1(n15889), .I2(n25059), .O(n25776) );
  INV1S U30046 ( .I(n25776), .O(n25778) );
  MOAI1S U30047 ( .A1(n25062), .A2(n25341), .B1(n25061), .B2(n25339), .O(
        n25063) );
  NR2 U30048 ( .I1(n15889), .I2(n25063), .O(n25834) );
  INV1S U30049 ( .I(n25834), .O(n25836) );
  MOAI1S U30050 ( .A1(n25341), .A2(n25066), .B1(n25339), .B2(n25065), .O(
        n25067) );
  NR2 U30051 ( .I1(n15889), .I2(n25067), .O(n25830) );
  ND2S U30052 ( .I1(n25830), .I2(gray_img[1895]), .O(n25069) );
  INV1S U30053 ( .I(gray_img[1895]), .O(n25070) );
  ND2S U30054 ( .I1(n27447), .I2(n25070), .O(n25068) );
  OAI112HS U30055 ( .C1(n25291), .C2(n25830), .A1(n25069), .B1(n25068), .O(
        n15487) );
  INV1S U30056 ( .I(gray_img[951]), .O(n25073) );
  ND2S U30057 ( .I1(n25070), .I2(n25848), .O(n25869) );
  INV1S U30058 ( .I(n25869), .O(n25071) );
  NR2 U30059 ( .I1(gray_img[2031]), .I2(gray_img[1903]), .O(n25868) );
  ND2S U30060 ( .I1(n25071), .I2(n25868), .O(n25072) );
  AOI22S U30061 ( .A1(n16006), .A2(n25073), .B1(n25315), .B2(n25072), .O(
        n25074) );
  ND2S U30062 ( .I1(n25291), .I2(n25074), .O(n25076) );
  AOI22S U30063 ( .A1(n25373), .A2(n25217), .B1(n25371), .B2(n25347), .O(
        n25075) );
  MUX2S U30064 ( .A(gray_img[951]), .B(n25076), .S(n26090), .O(n13814) );
  INV1S U30065 ( .I(gray_img[1663]), .O(n25077) );
  INV1S U30066 ( .I(gray_img[1791]), .O(n25995) );
  ND2S U30067 ( .I1(n25077), .I2(n25995), .O(n26017) );
  INV1S U30068 ( .I(n26017), .O(n25078) );
  NR2 U30069 ( .I1(gray_img[1783]), .I2(gray_img[1655]), .O(n26016) );
  ND2S U30070 ( .I1(n25078), .I2(n26016), .O(n25079) );
  AOI22S U30071 ( .A1(n16006), .A2(n25080), .B1(n25315), .B2(n25079), .O(
        n25081) );
  ND2S U30072 ( .I1(n25291), .I2(n25081), .O(n25083) );
  AOI22S U30073 ( .A1(n25103), .A2(n25283), .B1(n25356), .B2(n25282), .O(
        n25082) );
  MUX2S U30074 ( .A(gray_img[831]), .B(n25083), .S(n26073), .O(n13860) );
  NR2 U30075 ( .I1(gray_img[311]), .I2(gray_img[439]), .O(n26520) );
  INV1S U30076 ( .I(gray_img[447]), .O(n25084) );
  INV1S U30077 ( .I(gray_img[319]), .O(n26501) );
  ND2S U30078 ( .I1(n25084), .I2(n26501), .O(n26521) );
  AN2B1S U30079 ( .I1(n26520), .B1(n26521), .O(n25090) );
  AOI22S U30080 ( .A1(n25246), .A2(n25086), .B1(n25257), .B2(n25085), .O(
        n25087) );
  OA12S U30081 ( .B1(gray_img[159]), .B2(n29427), .A1(n27845), .O(n25088) );
  MOAI1S U30082 ( .A1(n27845), .A2(gray_img[159]), .B1(n25291), .B2(n25088), 
        .O(n25089) );
  OAI12HS U30083 ( .B1(n29680), .B2(n25090), .A1(n25089), .O(n13755) );
  INV1S U30084 ( .I(gray_img[1559]), .O(n25091) );
  INV1S U30085 ( .I(gray_img[1687]), .O(n26558) );
  ND2S U30086 ( .I1(n25091), .I2(n26558), .O(n26567) );
  INV1S U30087 ( .I(n26567), .O(n25092) );
  NR2 U30088 ( .I1(gray_img[1567]), .I2(gray_img[1695]), .O(n26566) );
  ND2S U30089 ( .I1(n25092), .I2(n26566), .O(n25093) );
  AOI22S U30090 ( .A1(n16006), .A2(n25094), .B1(n25315), .B2(n25093), .O(
        n25095) );
  ND2S U30091 ( .I1(n25291), .I2(n25095), .O(n25097) );
  AOI22S U30092 ( .A1(n25103), .A2(n25326), .B1(n25356), .B2(n25325), .O(
        n25096) );
  MUX2S U30093 ( .A(gray_img[783]), .B(n25097), .S(n29580), .O(n13896) );
  INV1S U30094 ( .I(gray_img[775]), .O(n25101) );
  INV1S U30095 ( .I(gray_img[1551]), .O(n25098) );
  ND2S U30096 ( .I1(n25098), .I2(n26587), .O(n26609) );
  INV1S U30097 ( .I(n26609), .O(n25099) );
  NR2 U30098 ( .I1(gray_img[1543]), .I2(gray_img[1671]), .O(n26608) );
  ND2S U30099 ( .I1(n25099), .I2(n26608), .O(n25100) );
  AOI22S U30100 ( .A1(n16006), .A2(n25101), .B1(n25315), .B2(n25100), .O(
        n25102) );
  ND2S U30101 ( .I1(n25291), .I2(n25102), .O(n25105) );
  AOI22S U30102 ( .A1(n25103), .A2(n25218), .B1(n25356), .B2(n25216), .O(
        n25104) );
  MUX2S U30103 ( .A(gray_img[775]), .B(n25105), .S(n29481), .O(n13902) );
  INV1S U30104 ( .I(gray_img[1031]), .O(n25106) );
  ND2S U30105 ( .I1(n25106), .I2(n26639), .O(n26648) );
  INV1S U30106 ( .I(n26648), .O(n25107) );
  NR2 U30107 ( .I1(gray_img[1039]), .I2(gray_img[1167]), .O(n26647) );
  ND2S U30108 ( .I1(n25107), .I2(n26647), .O(n25108) );
  AOI22S U30109 ( .A1(n16006), .A2(n29929), .B1(n25315), .B2(n25108), .O(
        n25109) );
  ND2S U30110 ( .I1(n25291), .I2(n25109), .O(n25111) );
  AOI22S U30111 ( .A1(n25218), .A2(n25195), .B1(n25216), .B2(n25333), .O(
        n25110) );
  MUX2S U30112 ( .A(gray_img[519]), .B(n25111), .S(n29740), .O(n14066) );
  ND2S U30113 ( .I1(n25112), .I2(n30114), .O(n25117) );
  AN2B1S U30114 ( .I1(n25114), .B1(n25113), .O(n25115) );
  OA22S U30115 ( .A1(gray_img[7]), .A2(n30005), .B1(n29680), .B2(n25115), .O(
        n25116) );
  OAI112HS U30116 ( .C1(n30114), .C2(n25118), .A1(n25117), .B1(n25116), .O(
        n13613) );
  MOAI1S U30117 ( .A1(n25254), .A2(n25341), .B1(n25271), .B2(n25339), .O(
        n25119) );
  NR2 U30118 ( .I1(n15889), .I2(n25119), .O(n27543) );
  INV1S U30119 ( .I(n27543), .O(n27545) );
  MOAI1S U30120 ( .A1(n25258), .A2(n25341), .B1(n25257), .B2(n25339), .O(
        n25121) );
  NR2 U30121 ( .I1(n15889), .I2(n25121), .O(n27388) );
  INV1S U30122 ( .I(n27388), .O(n27390) );
  INV1S U30123 ( .I(gray_img[55]), .O(n27734) );
  ND2S U30124 ( .I1(n25123), .I2(n27406), .O(n27429) );
  INV1S U30125 ( .I(n27429), .O(n25124) );
  NR2 U30126 ( .I1(gray_img[103]), .I2(gray_img[231]), .O(n27428) );
  ND2S U30127 ( .I1(n25124), .I2(n27428), .O(n25125) );
  AOI22S U30128 ( .A1(n16006), .A2(n27734), .B1(n25315), .B2(n25125), .O(
        n25126) );
  ND2S U30129 ( .I1(n25291), .I2(n25126), .O(n25128) );
  AOI22S U30130 ( .A1(n25373), .A2(n25273), .B1(n25371), .B2(n25271), .O(
        n25127) );
  MUX2S U30131 ( .A(gray_img[55]), .B(n25128), .S(n27550), .O(n14232) );
  MOAI1S U30132 ( .A1(n25367), .A2(n25341), .B1(n25370), .B2(n25339), .O(
        n25129) );
  NR2 U30133 ( .I1(n15889), .I2(n25129), .O(n27772) );
  INV1S U30134 ( .I(n27772), .O(n27774) );
  MOAI1S U30135 ( .A1(n25362), .A2(n25341), .B1(n25361), .B2(n25339), .O(
        n25131) );
  NR2 U30136 ( .I1(n15889), .I2(n25131), .O(n27446) );
  INV1S U30137 ( .I(n27446), .O(n27449) );
  INV1S U30138 ( .I(gray_img[1047]), .O(n25133) );
  INV1S U30139 ( .I(gray_img[1175]), .O(n29811) );
  ND2S U30140 ( .I1(n25133), .I2(n29811), .O(n29820) );
  INV1S U30141 ( .I(n29820), .O(n25134) );
  NR2 U30142 ( .I1(gray_img[1183]), .I2(gray_img[1055]), .O(n29819) );
  ND2S U30143 ( .I1(n25134), .I2(n29819), .O(n25135) );
  AOI22S U30144 ( .A1(n16006), .A2(n25136), .B1(n25315), .B2(n25135), .O(
        n25137) );
  ND2S U30145 ( .I1(n25291), .I2(n25137), .O(n25139) );
  AOI22S U30146 ( .A1(n25195), .A2(n25326), .B1(n25333), .B2(n25325), .O(
        n25138) );
  MUX2S U30147 ( .A(gray_img[527]), .B(n25139), .S(n29881), .O(n14057) );
  MOAI1S U30148 ( .A1(n25334), .A2(n25352), .B1(n25333), .B2(n25351), .O(
        n25140) );
  NR2 U30149 ( .I1(n15889), .I2(n25140), .O(n27103) );
  INV1S U30150 ( .I(n27103), .O(n27105) );
  MOAI1S U30151 ( .A1(n25342), .A2(n25352), .B1(n25340), .B2(n25351), .O(
        n25142) );
  NR2 U30152 ( .I1(n15889), .I2(n25142), .O(n26994) );
  INV1S U30153 ( .I(n26994), .O(n26996) );
  MUX2S U30154 ( .A(n27447), .B(n26994), .S(gray_img[735]), .O(n25143) );
  MOAI1S U30155 ( .A1(n25334), .A2(n25357), .B1(n25333), .B2(n25355), .O(
        n25144) );
  NR2 U30156 ( .I1(n15889), .I2(n25144), .O(n27011) );
  INV1S U30157 ( .I(n27011), .O(n27013) );
  MOAI1S U30158 ( .A1(n25342), .A2(n25357), .B1(n25340), .B2(n25355), .O(
        n25146) );
  NR2 U30159 ( .I1(n15889), .I2(n25146), .O(n27007) );
  INV1S U30160 ( .I(n27007), .O(n27009) );
  AN2B1S U30161 ( .I1(n25149), .B1(n25148), .O(n25153) );
  OA12S U30162 ( .B1(gray_img[431]), .B2(n29427), .A1(n25151), .O(n25150) );
  MOAI1S U30163 ( .A1(n25151), .A2(gray_img[431]), .B1(n25291), .B2(n25150), 
        .O(n25152) );
  OAI12HS U30164 ( .B1(n29680), .B2(n25153), .A1(n25152), .O(n14109) );
  MOAI1S U30165 ( .A1(n25342), .A2(n25366), .B1(n25340), .B2(n25365), .O(
        n25154) );
  NR2 U30166 ( .I1(n15889), .I2(n25154), .O(n27241) );
  INV1S U30167 ( .I(n27241), .O(n27243) );
  MOAI1S U30168 ( .A1(n25334), .A2(n25366), .B1(n25333), .B2(n25365), .O(
        n25156) );
  NR2 U30169 ( .I1(n15889), .I2(n25156), .O(n27131) );
  INV1S U30170 ( .I(n27131), .O(n27133) );
  INV1S U30171 ( .I(gray_img[591]), .O(n25158) );
  ND2S U30172 ( .I1(n25158), .I2(n27158), .O(n27167) );
  INV1S U30173 ( .I(n27167), .O(n25159) );
  NR2 U30174 ( .I1(gray_img[711]), .I2(gray_img[583]), .O(n27166) );
  ND2S U30175 ( .I1(n25159), .I2(n27166), .O(n25160) );
  AOI22S U30176 ( .A1(n16006), .A2(n27275), .B1(n25315), .B2(n25160), .O(
        n25161) );
  ND2S U30177 ( .I1(n25291), .I2(n25161), .O(n25164) );
  AOI22S U30178 ( .A1(n25162), .A2(n25194), .B1(n25361), .B2(n25193), .O(
        n25163) );
  MUX2S U30179 ( .A(gray_img[295]), .B(n25164), .S(n27252), .O(n14162) );
  MOAI1S U30180 ( .A1(n25348), .A2(n25366), .B1(n25347), .B2(n25365), .O(
        n25165) );
  NR2 U30181 ( .I1(n15889), .I2(n25165), .O(n27259) );
  INV1S U30182 ( .I(n27259), .O(n27261) );
  MOAI1S U30183 ( .A1(n25358), .A2(n25366), .B1(n25356), .B2(n25365), .O(
        n25167) );
  NR2 U30184 ( .I1(n15889), .I2(n25167), .O(n27188) );
  INV1S U30185 ( .I(n27188), .O(n27190) );
  MOAI1S U30186 ( .A1(n25357), .A2(n25301), .B1(n25355), .B2(n25300), .O(
        n25169) );
  NR2 U30187 ( .I1(n15889), .I2(n25169), .O(n28421) );
  INV1S U30188 ( .I(n28421), .O(n28423) );
  MOAI1S U30189 ( .A1(n25357), .A2(n25297), .B1(n25355), .B2(n25296), .O(
        n25171) );
  NR2 U30190 ( .I1(n15889), .I2(n25171), .O(n28269) );
  INV1S U30191 ( .I(n28269), .O(n28271) );
  MOAI1S U30192 ( .A1(n25352), .A2(n25297), .B1(n25351), .B2(n25296), .O(
        n25173) );
  NR2 U30193 ( .I1(n15889), .I2(n25173), .O(n28286) );
  INV1S U30194 ( .I(n28286), .O(n28288) );
  MOAI1S U30195 ( .A1(n25352), .A2(n25301), .B1(n25351), .B2(n25300), .O(
        n25175) );
  NR2 U30196 ( .I1(n15889), .I2(n25175), .O(n28282) );
  INV1S U30197 ( .I(n28282), .O(n28284) );
  MOAI1S U30198 ( .A1(n25357), .A2(n25287), .B1(n25355), .B2(n25286), .O(
        n25177) );
  NR2 U30199 ( .I1(n15889), .I2(n25177), .O(n28594) );
  INV1S U30200 ( .I(n28594), .O(n28596) );
  MOAI1S U30201 ( .A1(n25357), .A2(n25293), .B1(n25355), .B2(n25292), .O(
        n25179) );
  NR2 U30202 ( .I1(n15889), .I2(n25179), .O(n28340) );
  INV1S U30203 ( .I(n28340), .O(n28342) );
  MOAI1S U30204 ( .A1(n25352), .A2(n25287), .B1(n25351), .B2(n25286), .O(
        n25181) );
  NR2 U30205 ( .I1(n15889), .I2(n25181), .O(n28357) );
  INV1S U30206 ( .I(n28357), .O(n28359) );
  MOAI1S U30207 ( .A1(n25352), .A2(n25293), .B1(n25351), .B2(n25292), .O(
        n25183) );
  NR2 U30208 ( .I1(n15889), .I2(n25183), .O(n28353) );
  INV1S U30209 ( .I(n28353), .O(n28355) );
  MOAI1S U30210 ( .A1(n25366), .A2(n25297), .B1(n25365), .B2(n25296), .O(
        n25185) );
  NR2 U30211 ( .I1(n15889), .I2(n25185), .O(n28473) );
  INV1S U30212 ( .I(n28473), .O(n28475) );
  MOAI1S U30213 ( .A1(n25366), .A2(n25301), .B1(n25365), .B2(n25300), .O(
        n25187) );
  NR2 U30214 ( .I1(n15889), .I2(n25187), .O(n28478) );
  INV1S U30215 ( .I(n28478), .O(n28480) );
  INV1S U30216 ( .I(gray_img[1095]), .O(n25189) );
  INV1S U30217 ( .I(gray_img[1223]), .O(n28506) );
  ND2S U30218 ( .I1(n25189), .I2(n28506), .O(n28515) );
  INV1S U30219 ( .I(n28515), .O(n25190) );
  NR2 U30220 ( .I1(gray_img[1231]), .I2(gray_img[1103]), .O(n28514) );
  ND2S U30221 ( .I1(n25190), .I2(n28514), .O(n25191) );
  AOI22S U30222 ( .A1(n16006), .A2(n28632), .B1(n25315), .B2(n25191), .O(
        n25192) );
  ND2S U30223 ( .I1(n25291), .I2(n25192), .O(n25197) );
  AOI22S U30224 ( .A1(n25195), .A2(n25194), .B1(n25333), .B2(n25193), .O(
        n25196) );
  MUX2S U30225 ( .A(gray_img[551]), .B(n25197), .S(n28672), .O(n14030) );
  MOAI1S U30226 ( .A1(n25366), .A2(n25293), .B1(n25365), .B2(n25292), .O(
        n25198) );
  NR2 U30227 ( .I1(n15889), .I2(n25198), .O(n28558) );
  ND2S U30228 ( .I1(n28558), .I2(gray_img[1487]), .O(n25201) );
  OAI112HS U30229 ( .C1(n25291), .C2(n28558), .A1(n25201), .B1(n25200), .O(
        n15538) );
  MOAI1S U30230 ( .A1(n25366), .A2(n25287), .B1(n25365), .B2(n25286), .O(
        n25202) );
  NR2 U30231 ( .I1(n15889), .I2(n25202), .O(n28533) );
  ND2S U30232 ( .I1(n28533), .I2(gray_img[1359]), .O(n25205) );
  OAI112HS U30233 ( .C1(n25291), .C2(n28533), .A1(n25205), .B1(n25204), .O(
        n15554) );
  INV1S U30234 ( .I(n25206), .O(n25208) );
  ND2S U30235 ( .I1(n25208), .I2(n25207), .O(n25209) );
  AOI22S U30236 ( .A1(n16006), .A2(n25210), .B1(n25315), .B2(n25209), .O(
        n25211) );
  ND2S U30237 ( .I1(n25291), .I2(n25211), .O(n25212) );
  MUX2S U30238 ( .A(gray_img[679]), .B(n25212), .S(n28581), .O(n13944) );
  INV1S U30239 ( .I(gray_img[903]), .O(n29628) );
  INV1S U30240 ( .I(gray_img[1935]), .O(n29411) );
  INV1S U30241 ( .I(gray_img[1807]), .O(n29414) );
  ND2S U30242 ( .I1(n29411), .I2(n29414), .O(n29423) );
  INV1S U30243 ( .I(n29423), .O(n25213) );
  NR2 U30244 ( .I1(gray_img[1799]), .I2(gray_img[1927]), .O(n29422) );
  ND2S U30245 ( .I1(n25213), .I2(n29422), .O(n25214) );
  AOI22S U30246 ( .A1(n16006), .A2(n29628), .B1(n25315), .B2(n25214), .O(
        n25215) );
  ND2S U30247 ( .I1(n25291), .I2(n25215), .O(n25220) );
  AOI22S U30248 ( .A1(n25218), .A2(n25217), .B1(n25216), .B2(n25347), .O(
        n25219) );
  MUX2S U30249 ( .A(gray_img[903]), .B(n25220), .S(n30092), .O(n13838) );
  MOAI1S U30250 ( .A1(n25254), .A2(n25352), .B1(n25271), .B2(n25351), .O(
        n25221) );
  NR2 U30251 ( .I1(n15889), .I2(n25221), .O(n26707) );
  ND2S U30252 ( .I1(n26707), .I2(gray_img[95]), .O(n25224) );
  OAI112HS U30253 ( .C1(n25291), .C2(n26707), .A1(n25224), .B1(n25223), .O(
        n15656) );
  MOAI1S U30254 ( .A1(n25258), .A2(n25352), .B1(n25257), .B2(n25351), .O(
        n25225) );
  NR2 U30255 ( .I1(n15889), .I2(n25225), .O(n26724) );
  INV1S U30256 ( .I(n26724), .O(n26726) );
  MOAI1S U30257 ( .A1(n25258), .A2(n25357), .B1(n25257), .B2(n25355), .O(
        n25227) );
  NR2 U30258 ( .I1(n15889), .I2(n25227), .O(n26839) );
  INV1S U30259 ( .I(n26839), .O(n26841) );
  MOAI1S U30260 ( .A1(n25254), .A2(n25357), .B1(n25271), .B2(n25355), .O(
        n25229) );
  NR2 U30261 ( .I1(n15889), .I2(n25229), .O(n26720) );
  INV1S U30262 ( .I(n26720), .O(n26722) );
  MOAI1S U30263 ( .A1(n25362), .A2(n25357), .B1(n25361), .B2(n25355), .O(
        n25231) );
  NR2 U30264 ( .I1(n15889), .I2(n25231), .O(n26741) );
  INV1S U30265 ( .I(n26741), .O(n26743) );
  MOAI1S U30266 ( .A1(n25367), .A2(n25357), .B1(n25370), .B2(n25355), .O(
        n25233) );
  NR2 U30267 ( .I1(n15889), .I2(n25233), .O(n26745) );
  INV1S U30268 ( .I(n26745), .O(n26747) );
  MOAI1S U30269 ( .A1(n25367), .A2(n25352), .B1(n25370), .B2(n25351), .O(
        n25235) );
  NR2 U30270 ( .I1(n15889), .I2(n25235), .O(n27350) );
  INV1S U30271 ( .I(n27350), .O(n27352) );
  INV1S U30272 ( .I(gray_img[479]), .O(n26786) );
  MOAI1S U30273 ( .A1(n25362), .A2(n25352), .B1(n25361), .B2(n25351), .O(
        n25237) );
  NR2 U30274 ( .I1(n15889), .I2(n25237), .O(n26757) );
  INV1S U30275 ( .I(n26757), .O(n26759) );
  INV1S U30276 ( .I(gray_img[351]), .O(n25239) );
  INV1S U30277 ( .I(gray_img[175]), .O(n25242) );
  ND2S U30278 ( .I1(n25239), .I2(n26786), .O(n26795) );
  INV1S U30279 ( .I(n26795), .O(n25240) );
  NR2 U30280 ( .I1(gray_img[343]), .I2(gray_img[471]), .O(n26794) );
  ND2S U30281 ( .I1(n25240), .I2(n26794), .O(n25241) );
  AOI22S U30282 ( .A1(n16006), .A2(n25242), .B1(n25315), .B2(n25241), .O(
        n25243) );
  ND2S U30283 ( .I1(n25291), .I2(n25243), .O(n25248) );
  AOI22S U30284 ( .A1(n25246), .A2(n25245), .B1(n25257), .B2(n25244), .O(
        n25247) );
  MUX2S U30285 ( .A(gray_img[175]), .B(n25248), .S(n27356), .O(n14197) );
  AN2B1S U30286 ( .I1(n25250), .B1(n25249), .O(n25253) );
  OA12S U30287 ( .B1(gray_img[167]), .B2(n29427), .A1(n26932), .O(n25251) );
  MOAI1S U30288 ( .A1(n26932), .A2(gray_img[167]), .B1(n25291), .B2(n25251), 
        .O(n25252) );
  OAI12HS U30289 ( .B1(n29680), .B2(n25253), .A1(n25252), .O(n14206) );
  MOAI1S U30290 ( .A1(n25254), .A2(n25366), .B1(n25271), .B2(n25365), .O(
        n25255) );
  NR2 U30291 ( .I1(n15889), .I2(n25255), .O(n26877) );
  INV1S U30292 ( .I(n26877), .O(n26879) );
  MOAI1S U30293 ( .A1(n25258), .A2(n25366), .B1(n25257), .B2(n25365), .O(
        n25259) );
  NR2 U30294 ( .I1(n15889), .I2(n25259), .O(n26881) );
  INV1S U30295 ( .I(n26881), .O(n26883) );
  INV1S U30296 ( .I(gray_img[39]), .O(n25267) );
  INV1S U30297 ( .I(n25261), .O(n25263) );
  ND2S U30298 ( .I1(n25263), .I2(n25262), .O(n25264) );
  AOI22S U30299 ( .A1(n16006), .A2(n25267), .B1(n25315), .B2(n25264), .O(
        n25265) );
  ND2S U30300 ( .I1(n25291), .I2(n25265), .O(n25266) );
  MUX2S U30301 ( .A(gray_img[39]), .B(n25266), .S(n26924), .O(n14250) );
  INV1S U30302 ( .I(gray_img[23]), .O(n27863) );
  INV1S U30303 ( .I(gray_img[167]), .O(n26955) );
  ND2S U30304 ( .I1(n25267), .I2(n26955), .O(n26977) );
  INV1S U30305 ( .I(n26977), .O(n25268) );
  NR2 U30306 ( .I1(gray_img[47]), .I2(gray_img[175]), .O(n26976) );
  ND2S U30307 ( .I1(n25268), .I2(n26976), .O(n25269) );
  AOI22S U30308 ( .A1(n16006), .A2(n27863), .B1(n25315), .B2(n25269), .O(
        n25270) );
  ND2S U30309 ( .I1(n25291), .I2(n25270), .O(n25276) );
  AOI22S U30310 ( .A1(n25274), .A2(n25273), .B1(n25272), .B2(n25271), .O(
        n25275) );
  MUX2S U30311 ( .A(gray_img[23]), .B(n25276), .S(n27371), .O(n13795) );
  INV1S U30312 ( .I(gray_img[703]), .O(n25280) );
  INV1S U30313 ( .I(gray_img[1527]), .O(n25277) );
  ND2S U30314 ( .I1(n25277), .I2(n27917), .O(n27926) );
  INV1S U30315 ( .I(n27926), .O(n25278) );
  NR2 U30316 ( .I1(gray_img[1535]), .I2(gray_img[1407]), .O(n27925) );
  ND2S U30317 ( .I1(n25278), .I2(n27925), .O(n25279) );
  AOI22S U30318 ( .A1(n16006), .A2(n25280), .B1(n25315), .B2(n25279), .O(
        n25281) );
  ND2S U30319 ( .I1(n25291), .I2(n25281), .O(n25285) );
  AOI22S U30320 ( .A1(n25308), .A2(n25283), .B1(n25340), .B2(n25282), .O(
        n25284) );
  MUX2S U30321 ( .A(gray_img[703]), .B(n25285), .S(n28137), .O(n13924) );
  MOAI1S U30322 ( .A1(n25341), .A2(n25287), .B1(n25339), .B2(n25286), .O(
        n25288) );
  NR2 U30323 ( .I1(n15889), .I2(n25288), .O(n28201) );
  ND2S U30324 ( .I1(n28201), .I2(gray_img[1383]), .O(n25290) );
  INV1S U30325 ( .I(gray_img[1383]), .O(n28002) );
  OAI112HS U30326 ( .C1(n25291), .C2(n28201), .A1(n25290), .B1(n25289), .O(
        n15551) );
  MOAI1S U30327 ( .A1(n25341), .A2(n25293), .B1(n25339), .B2(n25292), .O(
        n25294) );
  NR2 U30328 ( .I1(n15889), .I2(n25294), .O(n27969) );
  INV1S U30329 ( .I(n27969), .O(n27971) );
  MOAI1S U30330 ( .A1(n25341), .A2(n25297), .B1(n25339), .B2(n25296), .O(
        n25298) );
  NR2 U30331 ( .I1(n15889), .I2(n25298), .O(n28029) );
  INV1S U30332 ( .I(n28029), .O(n28031) );
  MOAI1S U30333 ( .A1(n25341), .A2(n25301), .B1(n25339), .B2(n25300), .O(
        n25302) );
  NR2 U30334 ( .I1(n15889), .I2(n25302), .O(n28090) );
  INV1S U30335 ( .I(n28090), .O(n28092) );
  INV1S U30336 ( .I(gray_img[1431]), .O(n25304) );
  INV1S U30337 ( .I(gray_img[1303]), .O(n29759) );
  ND2S U30338 ( .I1(n25304), .I2(n29759), .O(n29781) );
  INV1S U30339 ( .I(n29781), .O(n25305) );
  NR2 U30340 ( .I1(gray_img[1311]), .I2(gray_img[1439]), .O(n29780) );
  ND2S U30341 ( .I1(n25305), .I2(n29780), .O(n25306) );
  AOI22S U30342 ( .A1(n16006), .A2(n29917), .B1(n25315), .B2(n25306), .O(
        n25307) );
  ND2S U30343 ( .I1(n25291), .I2(n25307), .O(n25310) );
  AOI22S U30344 ( .A1(n25326), .A2(n25308), .B1(n25325), .B2(n25340), .O(
        n25309) );
  MUX2S U30345 ( .A(gray_img[655]), .B(n25310), .S(n29898), .O(n13969) );
  INV1S U30346 ( .I(gray_img[671]), .O(n25316) );
  INV1S U30347 ( .I(n25311), .O(n25313) );
  ND2S U30348 ( .I1(n25313), .I2(n25312), .O(n25314) );
  AOI22S U30349 ( .A1(n16006), .A2(n25316), .B1(n25315), .B2(n25314), .O(
        n25317) );
  ND2S U30350 ( .I1(n25291), .I2(n25317), .O(n25318) );
  MUX2S U30351 ( .A(gray_img[671]), .B(n25318), .S(n29344), .O(n13952) );
  AN2B1S U30352 ( .I1(n25320), .B1(n25319), .O(n25323) );
  OA12S U30353 ( .B1(gray_img[135]), .B2(n29427), .A1(n30121), .O(n25321) );
  MOAI1S U30354 ( .A1(n30121), .A2(gray_img[135]), .B1(n25291), .B2(n25321), 
        .O(n25322) );
  OAI12HS U30355 ( .B1(n29680), .B2(n25323), .A1(n25322), .O(n13622) );
  NR2 U30356 ( .I1(gray_img[919]), .I2(gray_img[791]), .O(n29306) );
  INV1S U30357 ( .I(gray_img[799]), .O(n25324) );
  INV1S U30358 ( .I(gray_img[927]), .O(n29286) );
  ND2S U30359 ( .I1(n25324), .I2(n29286), .O(n29307) );
  AN2B1S U30360 ( .I1(n29306), .B1(n29307), .O(n25330) );
  AOI22S U30361 ( .A1(n25372), .A2(n25326), .B1(n25370), .B2(n25325), .O(
        n25327) );
  OA12S U30362 ( .B1(gray_img[399]), .B2(n29427), .A1(n30032), .O(n25328) );
  MOAI1S U30363 ( .A1(n30032), .A2(gray_img[399]), .B1(n25291), .B2(n25328), 
        .O(n25329) );
  OAI12HS U30364 ( .B1(n29680), .B2(n25330), .A1(n25329), .O(n15070) );
  MOAI1S U30365 ( .A1(n25358), .A2(n25341), .B1(n25356), .B2(n25339), .O(
        n25331) );
  NR2 U30366 ( .I1(n15889), .I2(n25331), .O(n26222) );
  INV1S U30367 ( .I(n26222), .O(n26224) );
  MOAI1S U30368 ( .A1(n25334), .A2(n25341), .B1(n25333), .B2(n25339), .O(
        n25335) );
  NR2 U30369 ( .I1(n15889), .I2(n25335), .O(n26158) );
  INV1S U30370 ( .I(n26158), .O(n26160) );
  MOAI1S U30371 ( .A1(n25348), .A2(n25341), .B1(n25347), .B2(n25339), .O(
        n25337) );
  NR2 U30372 ( .I1(n15889), .I2(n25337), .O(n27827) );
  INV1S U30373 ( .I(n27827), .O(n27829) );
  MOAI1S U30374 ( .A1(n25342), .A2(n25341), .B1(n25340), .B2(n25339), .O(
        n25343) );
  NR2 U30375 ( .I1(n15889), .I2(n25343), .O(n26153) );
  INV1S U30376 ( .I(n26153), .O(n26155) );
  MOAI1S U30377 ( .A1(n25348), .A2(n25357), .B1(n25347), .B2(n25355), .O(
        n25345) );
  NR2 U30378 ( .I1(n15889), .I2(n25345), .O(n27063) );
  INV1S U30379 ( .I(n27063), .O(n27065) );
  MOAI1S U30380 ( .A1(n25348), .A2(n25352), .B1(n25347), .B2(n25351), .O(
        n25349) );
  NR2 U30381 ( .I1(n15889), .I2(n25349), .O(n27079) );
  INV1S U30382 ( .I(n27079), .O(n27081) );
  MOAI1S U30383 ( .A1(n25358), .A2(n25352), .B1(n25356), .B2(n25351), .O(
        n25353) );
  NR2 U30384 ( .I1(n15889), .I2(n25353), .O(n30063) );
  INV1S U30385 ( .I(n30063), .O(n30065) );
  MOAI1S U30386 ( .A1(n25358), .A2(n25357), .B1(n25356), .B2(n25355), .O(
        n25359) );
  NR2 U30387 ( .I1(n15889), .I2(n25359), .O(n27067) );
  INV1S U30388 ( .I(n27067), .O(n27069) );
  MOAI1S U30389 ( .A1(n25362), .A2(n25366), .B1(n25361), .B2(n25365), .O(
        n25363) );
  NR2 U30390 ( .I1(n27447), .I2(n25363), .O(n26859) );
  INV1S U30391 ( .I(n26859), .O(n26861) );
  MOAI1S U30392 ( .A1(n25367), .A2(n25366), .B1(n25370), .B2(n25365), .O(
        n25368) );
  NR2 U30393 ( .I1(n15889), .I2(n25368), .O(n26940) );
  INV1S U30394 ( .I(n26940), .O(n26942) );
  NR2 U30395 ( .I1(gray_img[999]), .I2(gray_img[871]), .O(n26263) );
  INV1S U30396 ( .I(gray_img[1007]), .O(n26240) );
  INV1S U30397 ( .I(gray_img[879]), .O(n26243) );
  ND2S U30398 ( .I1(n26240), .I2(n26243), .O(n26264) );
  AN2B1S U30399 ( .I1(n26263), .B1(n26264), .O(n25378) );
  AOI22S U30400 ( .A1(n25373), .A2(n25372), .B1(n25371), .B2(n25370), .O(
        n25375) );
  OA12S U30401 ( .B1(gray_img[439]), .B2(n29427), .A1(n27834), .O(n25376) );
  MOAI1S U30402 ( .A1(n27834), .A2(gray_img[439]), .B1(n25291), .B2(n25376), 
        .O(n25377) );
  OAI12HS U30403 ( .B1(n29680), .B2(n25378), .A1(n25377), .O(n14100) );
  INV1S U30404 ( .I(n29825), .O(n25444) );
  INV1S U30405 ( .I(n29825), .O(n25448) );
  INV1S U30406 ( .I(n25651), .O(n25653) );
  MUX2S U30407 ( .A(n27447), .B(n25471), .S(gray_img[2014]), .O(n25381) );
  MUX2S U30408 ( .A(n27447), .B(n27011), .S(gray_img[598]), .O(n25385) );
  MUX2S U30409 ( .A(n27447), .B(n26724), .S(gray_img[222]), .O(n25386) );
  INV1S U30410 ( .I(n25647), .O(n25649) );
  MUX2S U30411 ( .A(n15889), .B(n27188), .S(gray_img[846]), .O(n25390) );
  MUX2S U30412 ( .A(n27447), .B(n28357), .S(gray_img[1374]), .O(n25392) );
  INV1S U30413 ( .I(n26707), .O(n26709) );
  MUX2S U30414 ( .A(n15889), .B(n27007), .S(gray_img[726]), .O(n25396) );
  MUX2S U30415 ( .A(n15889), .B(n27131), .S(gray_img[590]), .O(n25398) );
  MUX2S U30416 ( .A(n27447), .B(n26839), .S(gray_img[214]), .O(n25399) );
  MUX2S U30417 ( .A(n15889), .B(n28421), .S(gray_img[1110]), .O(n25400) );
  INV1S U30418 ( .I(n25475), .O(n25477) );
  ND2S U30419 ( .I1(n25759), .I2(gray_img[2006]), .O(n25405) );
  OAI112HS U30420 ( .C1(n29825), .C2(n25759), .A1(n25405), .B1(n25404), .O(
        n15278) );
  INV1S U30421 ( .I(n28558), .O(n28560) );
  MUX2S U30422 ( .A(n27447), .B(n28558), .S(gray_img[1486]), .O(n25406) );
  INV1S U30423 ( .I(n28533), .O(n28536) );
  MUX2S U30424 ( .A(n15889), .B(n28533), .S(gray_img[1358]), .O(n25407) );
  MUX2S U30425 ( .A(n27447), .B(n28340), .S(gray_img[1494]), .O(n25408) );
  MUX2S U30426 ( .A(n15889), .B(n27259), .S(gray_img[974]), .O(n25409) );
  MUX2S U30427 ( .A(n27447), .B(n26720), .S(gray_img[86]), .O(n25411) );
  MUX2S U30428 ( .A(n27447), .B(n30063), .S(gray_img[862]), .O(n25413) );
  MUX2S U30429 ( .A(n27447), .B(n28473), .S(gray_img[1230]), .O(n25416) );
  MUX2S U30430 ( .A(n27447), .B(n27103), .S(gray_img[606]), .O(n25418) );
  MUX2S U30431 ( .A(n15889), .B(n28282), .S(gray_img[1118]), .O(n25419) );
  MUX2S U30432 ( .A(n15889), .B(n27241), .S(gray_img[718]), .O(n25420) );
  MUX2S U30433 ( .A(n27447), .B(n27067), .S(gray_img[854]), .O(n25421) );
  INV1S U30434 ( .I(n25629), .O(n25631) );
  MUX2S U30435 ( .A(n27447), .B(n26757), .S(gray_img[350]), .O(n25426) );
  MUX2S U30436 ( .A(n15889), .B(n26940), .S(gray_img[462]), .O(n25427) );
  MUX2S U30437 ( .A(n15889), .B(n28286), .S(gray_img[1246]), .O(n25428) );
  MUX2S U30438 ( .A(n27447), .B(n25496), .S(gray_img[1750]), .O(n25429) );
  INV1S U30439 ( .I(n25830), .O(n25832) );
  MUX2S U30440 ( .A(n26158), .B(n15889), .S(n26200), .O(n25433) );
  MUX2S U30441 ( .A(n27447), .B(n27827), .S(gray_img[998]), .O(n25436) );
  INV1S U30442 ( .I(gray_img[742]), .O(n26199) );
  MUX2S U30443 ( .A(n26153), .B(n15889), .S(n26199), .O(n25437) );
  ND2S U30444 ( .I1(n28201), .I2(gray_img[1382]), .O(n25441) );
  INV1S U30445 ( .I(gray_img[1382]), .O(n27997) );
  OAI112HS U30446 ( .C1(n29825), .C2(n28201), .A1(n25441), .B1(n25440), .O(
        n15356) );
  MUX2S U30447 ( .A(n27447), .B(n25759), .S(gray_img[2005]), .O(n25449) );
  MUX2S U30448 ( .A(n27447), .B(n25759), .S(gray_img[2004]), .O(n25451) );
  MUX2S U30449 ( .A(n27447), .B(n25458), .S(gray_img[1875]), .O(n25452) );
  AO12S U30450 ( .B1(n15888), .B2(n25460), .A1(n25454), .O(n13849) );
  MUX2S U30451 ( .A(n27447), .B(n25458), .S(gray_img[1876]), .O(n25455) );
  MUX2S U30452 ( .A(n27447), .B(n25759), .S(gray_img[2002]), .O(n25457) );
  MUX2S U30453 ( .A(n28534), .B(n25759), .S(gray_img[2001]), .O(n25461) );
  MUX2S U30454 ( .A(n27447), .B(n25471), .S(gray_img[2010]), .O(n25465) );
  AO12S U30455 ( .B1(n15888), .B2(n25473), .A1(n25466), .O(n13818) );
  MUX2S U30456 ( .A(n27447), .B(n25475), .S(gray_img[1884]), .O(n25468) );
  MUX2S U30457 ( .A(n27447), .B(n25475), .S(gray_img[1883]), .O(n25469) );
  MUX2S U30458 ( .A(n28534), .B(n25475), .S(gray_img[1882]), .O(n25470) );
  MUX2S U30459 ( .A(n28534), .B(n25471), .S(gray_img[2009]), .O(n25472) );
  AO12S U30460 ( .B1(n15888), .B2(n25477), .A1(n25476), .O(n13848) );
  ND2S U30461 ( .I1(n15890), .I2(n25612), .O(n25478) );
  OAI112HS U30462 ( .C1(n25616), .C2(n25480), .A1(n25479), .B1(n25478), .O(
        n25481) );
  MUX2S U30463 ( .A(n27447), .B(n25492), .S(gray_img[1621]), .O(n25483) );
  MUX2S U30464 ( .A(n27447), .B(n25492), .S(gray_img[1620]), .O(n25484) );
  MUX2S U30465 ( .A(n27447), .B(n25492), .S(gray_img[1618]), .O(n25486) );
  MUX2S U30466 ( .A(n27447), .B(n25492), .S(gray_img[1617]), .O(n25487) );
  MUX2S U30467 ( .A(n27447), .B(n25496), .S(gray_img[1746]), .O(n25491) );
  MUX2S U30468 ( .A(n27447), .B(n25492), .S(gray_img[1616]), .O(n25493) );
  AO12S U30469 ( .B1(n15888), .B2(n25494), .A1(n25493), .O(n13913) );
  MUX2S U30470 ( .A(n27447), .B(n25496), .S(gray_img[1744]), .O(n25497) );
  AO12S U30471 ( .B1(n15888), .B2(n25498), .A1(n25497), .O(n13877) );
  MUX2S U30472 ( .A(n27447), .B(n25508), .S(gray_img[1756]), .O(n25500) );
  MUX2S U30473 ( .A(n27447), .B(n25508), .S(gray_img[1755]), .O(n25501) );
  AO12S U30474 ( .B1(n15888), .B2(n25510), .A1(n25503), .O(n13876) );
  MUX2S U30475 ( .A(n27447), .B(n25574), .S(gray_img[1629]), .O(n25504) );
  MUX2S U30476 ( .A(n27447), .B(n25574), .S(gray_img[1628]), .O(n25505) );
  MUX2S U30477 ( .A(n27447), .B(n25574), .S(gray_img[1626]), .O(n25507) );
  MUX2S U30478 ( .A(n27447), .B(n25508), .S(gray_img[1753]), .O(n25509) );
  FA1S U30479 ( .A(intadd_39_B_0_), .B(n25512), .CI(gray_img[1745]), .CO(
        n25513) );
  FA1S U30480 ( .A(gray_img[1746]), .B(n25514), .CI(n25513), .CO(n25515) );
  FA1S U30481 ( .A(gray_img[1747]), .B(n25516), .CI(n25515), .CO(n25517) );
  MXL2HS U30482 ( .A(gray_img[1622]), .B(gray_img[1750]), .S(n25538), .OB(
        n25553) );
  INV1S U30483 ( .I(gray_img[1630]), .O(n25535) );
  INV1S U30484 ( .I(gray_img[1629]), .O(n25533) );
  INV1S U30485 ( .I(gray_img[1628]), .O(n25531) );
  INV1S U30486 ( .I(gray_img[1627]), .O(n25529) );
  INV1S U30487 ( .I(gray_img[1626]), .O(n25527) );
  FA1S U30488 ( .A(gray_img[1753]), .B(gray_img[1752]), .CI(n25525), .CO(
        n25526) );
  MAO222S U30489 ( .A1(n25527), .B1(gray_img[1754]), .C1(n25526), .O(n25528)
         );
  FA1S U30490 ( .A(n25529), .B(gray_img[1755]), .CI(n25528), .CO(n25530) );
  FA1S U30491 ( .A(n25531), .B(gray_img[1756]), .CI(n25530), .CO(n25532) );
  MXL2HS U30492 ( .A(gray_img[1621]), .B(gray_img[1749]), .S(n25538), .OB(
        n25558) );
  MXL2HS U30493 ( .A(gray_img[1620]), .B(gray_img[1748]), .S(n25538), .OB(
        n25563) );
  MXL2HS U30494 ( .A(gray_img[1619]), .B(gray_img[1747]), .S(n25538), .OB(
        n25568) );
  MUX2S U30495 ( .A(gray_img[1626]), .B(gray_img[1754]), .S(n25577), .O(n25569) );
  MXL2HS U30496 ( .A(gray_img[1618]), .B(gray_img[1746]), .S(n25538), .OB(
        n25573) );
  MXL2HS U30497 ( .A(gray_img[1617]), .B(gray_img[1745]), .S(n25538), .OB(
        n25611) );
  MXL2HS U30498 ( .A(gray_img[1616]), .B(gray_img[1744]), .S(n25538), .OB(
        n25582) );
  MUX2S U30499 ( .A(gray_img[1625]), .B(gray_img[1753]), .S(n25577), .O(n25603) );
  OR2 U30500 ( .I1(n29680), .I2(n25547), .O(n25610) );
  INV1S U30501 ( .I(n25547), .O(n25548) );
  ND2S U30502 ( .I1(n25604), .I2(n25549), .O(n25552) );
  INV1S U30503 ( .I(n25605), .O(n25607) );
  MUX2S U30504 ( .A(n25928), .B(n25605), .S(gray_img[814]), .O(n25550) );
  OA12S U30505 ( .B1(n29825), .B2(n25607), .A1(n25550), .O(n25551) );
  OAI112HS U30506 ( .C1(n25553), .C2(n25610), .A1(n25552), .B1(n25551), .O(
        n13873) );
  ND2S U30507 ( .I1(n25604), .I2(n25554), .O(n25557) );
  MUX2S U30508 ( .A(n25928), .B(n25605), .S(gray_img[813]), .O(n25555) );
  OAI112HS U30509 ( .C1(n25558), .C2(n25610), .A1(n25557), .B1(n25556), .O(
        n13874) );
  ND2S U30510 ( .I1(n25604), .I2(n25559), .O(n25562) );
  MUX2S U30511 ( .A(n25928), .B(n25605), .S(gray_img[812]), .O(n25560) );
  OA12S U30512 ( .B1(n29837), .B2(n25607), .A1(n25560), .O(n25561) );
  OAI112HS U30513 ( .C1(n25563), .C2(n25610), .A1(n25562), .B1(n25561), .O(
        n13875) );
  ND2S U30514 ( .I1(n25604), .I2(n25564), .O(n25567) );
  OAI112HS U30515 ( .C1(n25568), .C2(n25610), .A1(n25567), .B1(n25566), .O(
        n13645) );
  ND2S U30516 ( .I1(n25604), .I2(n25569), .O(n25572) );
  OAI112HS U30517 ( .C1(n25573), .C2(n25610), .A1(n25572), .B1(n25571), .O(
        n13666) );
  AO12S U30518 ( .B1(n15888), .B2(n25576), .A1(n25575), .O(n13912) );
  MUX2S U30519 ( .A(gray_img[1624]), .B(gray_img[1752]), .S(n25577), .O(n25578) );
  ND2S U30520 ( .I1(n25604), .I2(n25578), .O(n25581) );
  MUX2S U30521 ( .A(n25928), .B(n25605), .S(gray_img[808]), .O(n25579) );
  OAI112HS U30522 ( .C1(n25582), .C2(n25610), .A1(n25581), .B1(n25580), .O(
        n13717) );
  ND2S U30523 ( .I1(n15891), .I2(n25612), .O(n25583) );
  OAI112HS U30524 ( .C1(n25616), .C2(n25585), .A1(n25584), .B1(n25583), .O(
        n25586) );
  OAI112HS U30525 ( .C1(n25616), .C2(n25590), .A1(n25589), .B1(n25588), .O(
        n25591) );
  OAI112HS U30526 ( .C1(n25616), .C2(n25595), .A1(n25594), .B1(n25593), .O(
        n25596) );
  OAI112HS U30527 ( .C1(n25616), .C2(n25600), .A1(n25599), .B1(n25598), .O(
        n25601) );
  ND2S U30528 ( .I1(n25604), .I2(n25603), .O(n25609) );
  OAI112HS U30529 ( .C1(n25611), .C2(n25610), .A1(n25609), .B1(n25608), .O(
        n13690) );
  OAI112HS U30530 ( .C1(n25616), .C2(n25615), .A1(n25614), .B1(n25613), .O(
        n25617) );
  MUX2S U30531 ( .A(n27447), .B(n25629), .S(gray_img[1869]), .O(n25620) );
  AO12S U30532 ( .B1(n15888), .B2(n25631), .A1(n25624), .O(n13850) );
  MUX2S U30533 ( .A(n27447), .B(n28801), .S(gray_img[1997]), .O(n25625) );
  MUX2S U30534 ( .A(n27447), .B(n28801), .S(gray_img[1994]), .O(n25628) );
  MUX2S U30535 ( .A(n27447), .B(n28801), .S(gray_img[1993]), .O(n25632) );
  OAI112HS U30536 ( .C1(n25755), .C2(n25635), .A1(n25634), .B1(n25633), .O(
        n25636) );
  MUX2S U30537 ( .A(n27447), .B(n25647), .S(gray_img[1741]), .O(n25638) );
  AO12S U30538 ( .B1(n15888), .B2(n25649), .A1(n25642), .O(n13882) );
  MUX2S U30539 ( .A(n27447), .B(n25651), .S(gray_img[1612]), .O(n25644) );
  MUX2S U30540 ( .A(n15889), .B(n25651), .S(gray_img[1611]), .O(n25645) );
  MUX2S U30541 ( .A(n27447), .B(n25651), .S(gray_img[1610]), .O(n25646) );
  MUX2S U30542 ( .A(n27447), .B(n25651), .S(gray_img[1609]), .O(n25650) );
  AO12S U30543 ( .B1(n15888), .B2(n25653), .A1(n25652), .O(n13914) );
  INV1S U30544 ( .I(gray_img[1607]), .O(n25678) );
  INV1S U30545 ( .I(gray_img[1605]), .O(n25674) );
  INV1S U30546 ( .I(gray_img[1602]), .O(n25668) );
  FA1S U30547 ( .A(gray_img[1729]), .B(gray_img[1728]), .CI(intadd_42_CI), 
        .CO(n25667) );
  FA1S U30548 ( .A(n25668), .B(gray_img[1730]), .CI(n25667), .CO(n25669) );
  FA1S U30549 ( .A(n25670), .B(gray_img[1731]), .CI(n25669), .CO(n25671) );
  FA1S U30550 ( .A(n25672), .B(gray_img[1732]), .CI(n25671), .CO(n25673) );
  MXL2HS U30551 ( .A(gray_img[1606]), .B(gray_img[1734]), .S(n25741), .OB(
        n25692) );
  MXL2HS U30552 ( .A(gray_img[1605]), .B(gray_img[1733]), .S(n25741), .OB(
        n25697) );
  MXL2HS U30553 ( .A(gray_img[1604]), .B(gray_img[1732]), .S(n25741), .OB(
        n25702) );
  MXL2HS U30554 ( .A(gray_img[1603]), .B(gray_img[1731]), .S(n25741), .OB(
        n25707) );
  MXL2HS U30555 ( .A(gray_img[1602]), .B(gray_img[1730]), .S(n25741), .OB(
        n25712) );
  MXL2HS U30556 ( .A(gray_img[1601]), .B(gray_img[1729]), .S(n25741), .OB(
        n25717) );
  INV1S U30557 ( .I(n25689), .O(n25688) );
  NR2 U30558 ( .I1(n29680), .I2(n25688), .O(n25750) );
  ND2S U30559 ( .I1(n15890), .I2(n25744), .O(n25690) );
  OAI112HS U30560 ( .C1(n25740), .C2(n25692), .A1(n25691), .B1(n25690), .O(
        n25693) );
  OAI112HS U30561 ( .C1(n25740), .C2(n25697), .A1(n25696), .B1(n25695), .O(
        n25698) );
  OAI112HS U30562 ( .C1(n25740), .C2(n25702), .A1(n25701), .B1(n25700), .O(
        n25703) );
  OAI112HS U30563 ( .C1(n25740), .C2(n25707), .A1(n25706), .B1(n25705), .O(
        n25708) );
  OAI112HS U30564 ( .C1(n25740), .C2(n25712), .A1(n25711), .B1(n25710), .O(
        n25713) );
  OAI112HS U30565 ( .C1(n25740), .C2(n25717), .A1(n25716), .B1(n25715), .O(
        n25718) );
  OAI112HS U30566 ( .C1(n25755), .C2(n25722), .A1(n25721), .B1(n25720), .O(
        n25723) );
  OAI112HS U30567 ( .C1(n25755), .C2(n25727), .A1(n25726), .B1(n25725), .O(
        n25728) );
  OAI112HS U30568 ( .C1(n25755), .C2(n25732), .A1(n25731), .B1(n25730), .O(
        n25733) );
  OAI112HS U30569 ( .C1(n25755), .C2(n25737), .A1(n25736), .B1(n25735), .O(
        n25738) );
  INV1S U30570 ( .I(n25740), .O(n25743) );
  MUX2S U30571 ( .A(gray_img[1600]), .B(gray_img[1728]), .S(n25741), .O(n25742) );
  ND2S U30572 ( .I1(n25743), .I2(n25742), .O(n25747) );
  ND2S U30573 ( .I1(n15888), .I2(n25744), .O(n25745) );
  ND3S U30574 ( .I1(n25747), .I2(n25746), .I3(n25745), .O(n25748) );
  OAI112HS U30575 ( .C1(n25755), .C2(n25754), .A1(n25753), .B1(n25752), .O(
        n25756) );
  AO12S U30576 ( .B1(n15888), .B2(n25761), .A1(n25760), .O(n13819) );
  OA12S U30577 ( .B1(n29825), .B2(n28809), .A1(n25763), .O(n25764) );
  OAI112HS U30578 ( .C1(n25766), .C2(n28812), .A1(n25765), .B1(n25764), .O(
        n13617) );
  MUX2S U30579 ( .A(n27447), .B(n25776), .S(gray_img[1764]), .O(n25768) );
  MUX2S U30580 ( .A(n27447), .B(n25776), .S(gray_img[1760]), .O(n25771) );
  AO12S U30581 ( .B1(n15888), .B2(n25778), .A1(n25771), .O(n13871) );
  MUX2S U30582 ( .A(n27447), .B(n25897), .S(gray_img[1637]), .O(n25772) );
  MUX2S U30583 ( .A(n27447), .B(n25776), .S(gray_img[1761]), .O(n25777) );
  MUX2S U30584 ( .A(n27447), .B(n25897), .S(gray_img[1633]), .O(n25779) );
  INV1S U30585 ( .I(gray_img[1643]), .O(n25784) );
  INV1S U30586 ( .I(gray_img[1641]), .O(n25780) );
  INV1S U30587 ( .I(gray_img[1638]), .O(n25802) );
  INV1S U30588 ( .I(gray_img[1637]), .O(n25800) );
  INV1S U30589 ( .I(gray_img[1636]), .O(n25798) );
  INV1S U30590 ( .I(gray_img[1635]), .O(n25796) );
  MAO222S U30591 ( .A1(gray_img[1761]), .B1(gray_img[1760]), .C1(intadd_36_CI), 
        .O(n25793) );
  FA1S U30592 ( .A(n25794), .B(gray_img[1762]), .CI(n25793), .CO(n25795) );
  FA1S U30593 ( .A(n25796), .B(gray_img[1763]), .CI(n25795), .CO(n25797) );
  FA1S U30594 ( .A(n25798), .B(gray_img[1764]), .CI(n25797), .CO(n25799) );
  MXL2HS U30595 ( .A(gray_img[1638]), .B(gray_img[1766]), .S(n25900), .OB(
        n25818) );
  MXL2HS U30596 ( .A(gray_img[1637]), .B(gray_img[1765]), .S(n25900), .OB(
        n25879) );
  MXL2HS U30597 ( .A(gray_img[1636]), .B(gray_img[1764]), .S(n25900), .OB(
        n25884) );
  MXL2HS U30598 ( .A(gray_img[1635]), .B(gray_img[1763]), .S(n25900), .OB(
        n25889) );
  MXL2HS U30599 ( .A(gray_img[1634]), .B(gray_img[1762]), .S(n25900), .OB(
        n25894) );
  MUX2S U30600 ( .A(gray_img[1641]), .B(gray_img[1769]), .S(n25805), .O(n25935) );
  MXL2HS U30601 ( .A(gray_img[1633]), .B(gray_img[1761]), .S(n25900), .OB(
        n25932) );
  INV1S U30602 ( .I(n25815), .O(n25814) );
  NR2 U30603 ( .I1(n29680), .I2(n25814), .O(n25936) );
  ND2S U30604 ( .I1(n15890), .I2(n25929), .O(n25816) );
  OAI112HS U30605 ( .C1(n25933), .C2(n25818), .A1(n25817), .B1(n25816), .O(
        n25819) );
  MUX2S U30606 ( .A(n27447), .B(n25830), .S(gray_img[1890]), .O(n25824) );
  MUX2S U30607 ( .A(n27447), .B(n25834), .S(gray_img[2018]), .O(n25829) );
  AO12S U30608 ( .B1(n19092), .B2(n25832), .A1(n25831), .O(n13847) );
  MUX2S U30609 ( .A(n27447), .B(n25834), .S(gray_img[2017]), .O(n25833) );
  AO12S U30610 ( .B1(n15888), .B2(n25836), .A1(n25835), .O(n13816) );
  FA1S U30611 ( .A(gray_img[1888]), .B(gray_img[1889]), .CI(intadd_4_CI), .CO(
        n25837) );
  FA1S U30612 ( .A(n25838), .B(gray_img[1890]), .CI(n25837), .CO(n25839) );
  FA1S U30613 ( .A(n25840), .B(gray_img[1891]), .CI(n25839), .CO(n25841) );
  FA1S U30614 ( .A(intadd_5_B_0_), .B(gray_img[1897]), .CI(intadd_5_CI), .CO(
        n25849) );
  FA1S U30615 ( .A(n25850), .B(gray_img[1898]), .CI(n25849), .CO(n25851) );
  FA1S U30616 ( .A(n25852), .B(gray_img[1899]), .CI(n25851), .CO(n25853) );
  MXL2HS U30617 ( .A(gray_img[2030]), .B(gray_img[1902]), .S(n26087), .OB(
        n25874) );
  MXL2HS U30618 ( .A(gray_img[2029]), .B(gray_img[1901]), .S(n26087), .OB(
        n25910) );
  MXL2HS U30619 ( .A(gray_img[2028]), .B(gray_img[1900]), .S(n26087), .OB(
        n25915) );
  MXL2HS U30620 ( .A(gray_img[2027]), .B(gray_img[1899]), .S(n26087), .OB(
        n25920) );
  MXL2HS U30621 ( .A(gray_img[2026]), .B(gray_img[1898]), .S(n26087), .OB(
        n25925) );
  MXL2HS U30622 ( .A(gray_img[2025]), .B(gray_img[1897]), .S(n26087), .OB(
        n25939) );
  INV1S U30623 ( .I(n25871), .O(n25870) );
  NR2 U30624 ( .I1(n29680), .I2(n25870), .O(n26096) );
  OR2 U30625 ( .I1(n29680), .I2(n25871), .O(n26086) );
  OAI112HS U30626 ( .C1(n26086), .C2(n25874), .A1(n25873), .B1(n25872), .O(
        n25875) );
  ND2S U30627 ( .I1(n15891), .I2(n25929), .O(n25877) );
  OAI112HS U30628 ( .C1(n25933), .C2(n25879), .A1(n25878), .B1(n25877), .O(
        n25880) );
  OAI112HS U30629 ( .C1(n25933), .C2(n25884), .A1(n25883), .B1(n25882), .O(
        n25885) );
  ND2S U30630 ( .I1(n15927), .I2(n25929), .O(n25887) );
  OAI112HS U30631 ( .C1(n25933), .C2(n25889), .A1(n25888), .B1(n25887), .O(
        n25890) );
  ND2S U30632 ( .I1(n15934), .I2(n25929), .O(n25892) );
  OAI112HS U30633 ( .C1(n25933), .C2(n25894), .A1(n25893), .B1(n25892), .O(
        n25895) );
  AO12S U30634 ( .B1(n15888), .B2(n25899), .A1(n25898), .O(n13911) );
  INV1S U30635 ( .I(n25933), .O(n25902) );
  MUX2S U30636 ( .A(gray_img[1632]), .B(gray_img[1760]), .S(n25900), .O(n25901) );
  ND2S U30637 ( .I1(n25902), .I2(n25901), .O(n25905) );
  ND2S U30638 ( .I1(n15888), .I2(n25929), .O(n25903) );
  OAI112HS U30639 ( .C1(n26086), .C2(n25910), .A1(n25909), .B1(n25908), .O(
        n25911) );
  OAI112HS U30640 ( .C1(n26086), .C2(n25915), .A1(n25914), .B1(n25913), .O(
        n25916) );
  OAI112HS U30641 ( .C1(n26086), .C2(n25920), .A1(n25919), .B1(n25918), .O(
        n25921) );
  OAI112HS U30642 ( .C1(n26086), .C2(n25925), .A1(n25924), .B1(n25923), .O(
        n25926) );
  ND2S U30643 ( .I1(n15928), .I2(n25929), .O(n25930) );
  OAI112HS U30644 ( .C1(n25933), .C2(n25932), .A1(n25931), .B1(n25930), .O(
        n25934) );
  OAI112HS U30645 ( .C1(n26086), .C2(n25939), .A1(n25938), .B1(n25937), .O(
        n25940) );
  ND2S U30646 ( .I1(n29837), .I2(n25942), .O(n25945) );
  INV1S U30647 ( .I(gray_img[2036]), .O(n25963) );
  ND2S U30648 ( .I1(n25943), .I2(n25963), .O(n25944) );
  MOAI1S U30649 ( .A1(gray_img[2036]), .A2(n30005), .B1(n25945), .B2(n25944), 
        .O(n14878) );
  INV1S U30650 ( .I(gray_img[2047]), .O(n25957) );
  INV1S U30651 ( .I(gray_img[2046]), .O(n25955) );
  INV1S U30652 ( .I(gray_img[2045]), .O(n25953) );
  INV1S U30653 ( .I(gray_img[2044]), .O(n25951) );
  INV1S U30654 ( .I(gray_img[2043]), .O(n25949) );
  FA1S U30655 ( .A(gray_img[1912]), .B(intadd_2_A_0_), .CI(gray_img[1913]), 
        .CO(n25946) );
  FA1S U30656 ( .A(gray_img[1914]), .B(n25947), .CI(n25946), .CO(n25948) );
  FA1S U30657 ( .A(gray_img[1915]), .B(n25949), .CI(n25948), .CO(n25950) );
  FA1S U30658 ( .A(gray_img[1916]), .B(n25951), .CI(n25950), .CO(n25952) );
  FA1S U30659 ( .A(gray_img[1917]), .B(n25953), .CI(n25952), .CO(n25954) );
  MXL2HS U30660 ( .A(gray_img[2046]), .B(gray_img[1918]), .S(n28715), .OB(
        n25981) );
  INV1S U30661 ( .I(gray_img[2038]), .O(n25967) );
  INV1S U30662 ( .I(gray_img[2037]), .O(n25965) );
  INV1S U30663 ( .I(gray_img[2035]), .O(n25961) );
  INV1S U30664 ( .I(gray_img[2034]), .O(n25959) );
  FA1S U30665 ( .A(gray_img[1905]), .B(gray_img[1904]), .CI(intadd_1_CI), .CO(
        n25958) );
  MXL2HS U30666 ( .A(gray_img[2045]), .B(gray_img[1917]), .S(n28715), .OB(
        n26055) );
  MXL2HS U30667 ( .A(gray_img[2044]), .B(gray_img[1916]), .S(n28715), .OB(
        n26060) );
  MXL2HS U30668 ( .A(gray_img[2043]), .B(gray_img[1915]), .S(n28715), .OB(
        n26065) );
  MXL2HS U30669 ( .A(gray_img[2042]), .B(gray_img[1914]), .S(n28715), .OB(
        n26070) );
  MXL2HS U30670 ( .A(gray_img[2041]), .B(gray_img[1913]), .S(n28715), .OB(
        n26083) );
  MUX2S U30671 ( .A(gray_img[2032]), .B(gray_img[1904]), .S(n25970), .O(n28723) );
  FA1S U30672 ( .A(n26085), .B(n26083), .CI(n28723), .CO(n25971) );
  INV1S U30673 ( .I(n25978), .O(n25977) );
  NR2 U30674 ( .I1(n29680), .I2(n25977), .O(n28724) );
  OR2 U30675 ( .I1(n29680), .I2(n25978), .O(n28714) );
  ND2S U30676 ( .I1(n15890), .I2(n28718), .O(n25979) );
  OAI112HS U30677 ( .C1(n28714), .C2(n25981), .A1(n25980), .B1(n25979), .O(
        n25982) );
  INV1S U30678 ( .I(gray_img[1790]), .O(n25993) );
  INV1S U30679 ( .I(gray_img[1789]), .O(n25991) );
  INV1S U30680 ( .I(gray_img[1788]), .O(n25989) );
  INV1S U30681 ( .I(gray_img[1786]), .O(n25985) );
  MAO222S U30682 ( .A1(gray_img[1657]), .B1(gray_img[1656]), .C1(intadd_32_CI), 
        .O(n25984) );
  FA1S U30683 ( .A(n25985), .B(gray_img[1658]), .CI(n25984), .CO(n25986) );
  FA1S U30684 ( .A(n25987), .B(gray_img[1659]), .CI(n25986), .CO(n25988) );
  FA1S U30685 ( .A(n25989), .B(gray_img[1660]), .CI(n25988), .CO(n25990) );
  INV1S U30686 ( .I(gray_img[1783]), .O(n26008) );
  INV1S U30687 ( .I(gray_img[1782]), .O(n26006) );
  INV1S U30688 ( .I(gray_img[1781]), .O(n26004) );
  INV1S U30689 ( .I(gray_img[1778]), .O(n25998) );
  MXL2HS U30690 ( .A(gray_img[1782]), .B(gray_img[1654]), .S(n26045), .OB(
        n26022) );
  MXL2HS U30691 ( .A(gray_img[1781]), .B(gray_img[1653]), .S(n26045), .OB(
        n26027) );
  MXL2HS U30692 ( .A(gray_img[1780]), .B(gray_img[1652]), .S(n26045), .OB(
        n26032) );
  MXL2HS U30693 ( .A(gray_img[1779]), .B(gray_img[1651]), .S(n26045), .OB(
        n26037) );
  MXL2HS U30694 ( .A(gray_img[1778]), .B(gray_img[1650]), .S(n26045), .OB(
        n26042) );
  MXL2HS U30695 ( .A(gray_img[1777]), .B(gray_img[1649]), .S(n26045), .OB(
        n26076) );
  INV1S U30696 ( .I(n26019), .O(n26018) );
  NR2 U30697 ( .I1(n29680), .I2(n26018), .O(n26080) );
  ND2S U30698 ( .I1(n15890), .I2(n26073), .O(n26020) );
  OAI112HS U30699 ( .C1(n26077), .C2(n26022), .A1(n26021), .B1(n26020), .O(
        n26023) );
  OAI112HS U30700 ( .C1(n26077), .C2(n26027), .A1(n26026), .B1(n26025), .O(
        n26028) );
  OAI112HS U30701 ( .C1(n26077), .C2(n26032), .A1(n26031), .B1(n26030), .O(
        n26033) );
  OAI112HS U30702 ( .C1(n26077), .C2(n26037), .A1(n26036), .B1(n26035), .O(
        n26038) );
  OAI112HS U30703 ( .C1(n26077), .C2(n26042), .A1(n26041), .B1(n26040), .O(
        n26043) );
  INV1S U30704 ( .I(n26077), .O(n26047) );
  MUX2S U30705 ( .A(gray_img[1776]), .B(gray_img[1648]), .S(n26045), .O(n26046) );
  ND2S U30706 ( .I1(n26047), .I2(n26046), .O(n26050) );
  ND2S U30707 ( .I1(n15888), .I2(n26073), .O(n26048) );
  ND3S U30708 ( .I1(n26050), .I2(n26049), .I3(n26048), .O(n26051) );
  ND2S U30709 ( .I1(n15891), .I2(n28718), .O(n26053) );
  OAI112HS U30710 ( .C1(n28714), .C2(n26055), .A1(n26054), .B1(n26053), .O(
        n26056) );
  OAI112HS U30711 ( .C1(n28714), .C2(n26060), .A1(n26059), .B1(n26058), .O(
        n26061) );
  OAI112HS U30712 ( .C1(n28714), .C2(n26065), .A1(n26064), .B1(n26063), .O(
        n26066) );
  OAI112HS U30713 ( .C1(n28714), .C2(n26070), .A1(n26069), .B1(n26068), .O(
        n26071) );
  OAI112HS U30714 ( .C1(n26077), .C2(n26076), .A1(n26075), .B1(n26074), .O(
        n26078) );
  OAI112HS U30715 ( .C1(n28714), .C2(n26083), .A1(n26082), .B1(n26081), .O(
        n26084) );
  INV1S U30716 ( .I(n26086), .O(n26089) );
  MUX2S U30717 ( .A(gray_img[2024]), .B(gray_img[1896]), .S(n26087), .O(n26088) );
  ND2S U30718 ( .I1(n26089), .I2(n26088), .O(n26093) );
  ND2S U30719 ( .I1(n15888), .I2(n26090), .O(n26091) );
  ND3S U30720 ( .I1(n26093), .I2(n26092), .I3(n26091), .O(n26094) );
  INV1S U30721 ( .I(gray_img[819]), .O(n26102) );
  FA1S U30722 ( .A(n26098), .B(n26097), .CI(gray_img[945]), .CO(n26099) );
  FA1S U30723 ( .A(gray_img[946]), .B(n26100), .CI(n26099), .CO(n26101) );
  FA1S U30724 ( .A(gray_img[947]), .B(n26102), .CI(n26101), .CO(n26103) );
  MXL2HS U30725 ( .A(gray_img[822]), .B(gray_img[950]), .S(n26124), .OB(n26139) );
  INV1S U30726 ( .I(gray_img[957]), .O(n26119) );
  INV1S U30727 ( .I(gray_img[956]), .O(n26117) );
  INV1S U30728 ( .I(gray_img[955]), .O(n26115) );
  INV1S U30729 ( .I(gray_img[953]), .O(n26111) );
  FA1S U30730 ( .A(gray_img[825]), .B(gray_img[824]), .CI(n26111), .CO(n26112)
         );
  FA1S U30731 ( .A(n26113), .B(gray_img[826]), .CI(n26112), .CO(n26114) );
  FA1S U30732 ( .A(n26115), .B(gray_img[827]), .CI(n26114), .CO(n26116) );
  FA1S U30733 ( .A(n26117), .B(gray_img[828]), .CI(n26116), .CO(n26118) );
  MXL2HS U30734 ( .A(gray_img[821]), .B(gray_img[949]), .S(n26124), .OB(n28259) );
  MXL2HS U30735 ( .A(gray_img[820]), .B(gray_img[948]), .S(n26124), .OB(n28225) );
  MXL2HS U30736 ( .A(gray_img[819]), .B(gray_img[947]), .S(n26124), .OB(n28230) );
  MXL2HS U30737 ( .A(gray_img[818]), .B(gray_img[946]), .S(n26124), .OB(n28235) );
  MXL2HS U30738 ( .A(gray_img[816]), .B(gray_img[944]), .S(n26124), .OB(n28734) );
  MXL2HS U30739 ( .A(gray_img[817]), .B(gray_img[945]), .S(n26124), .OB(n28245) );
  OA12S U30740 ( .B1(gray_img[414]), .B2(n29427), .A1(n28728), .O(n26136) );
  MOAI1S U30741 ( .A1(n28728), .A2(gray_img[414]), .B1(n29825), .B2(n26136), 
        .O(n26137) );
  OAI112HS U30742 ( .C1(n26139), .C2(n28733), .A1(n26138), .B1(n26137), .O(
        n15271) );
  OA12S U30743 ( .B1(n29825), .B2(n29046), .A1(n26141), .O(n26142) );
  OAI112HS U30744 ( .C1(n26144), .C2(n29049), .A1(n26143), .B1(n26142), .O(
        n14049) );
  MUX2S U30745 ( .A(n15889), .B(n26153), .S(gray_img[741]), .O(n26145) );
  MUX2S U30746 ( .A(n27447), .B(n26153), .S(gray_img[739]), .O(n26147) );
  MUX2S U30747 ( .A(n15889), .B(n26153), .S(gray_img[738]), .O(n26148) );
  MUX2S U30748 ( .A(n15889), .B(n26153), .S(gray_img[736]), .O(n26149) );
  AO12S U30749 ( .B1(n15888), .B2(n26155), .A1(n26149), .O(n14152) );
  MUX2S U30750 ( .A(n15889), .B(n26158), .S(gray_img[612]), .O(n26150) );
  MUX2S U30751 ( .A(n15889), .B(n26158), .S(gray_img[611]), .O(n26151) );
  MUX2S U30752 ( .A(n27447), .B(n26158), .S(gray_img[610]), .O(n26152) );
  MUX2S U30753 ( .A(n15889), .B(n26158), .S(gray_img[609]), .O(n26156) );
  MUX2S U30754 ( .A(n27447), .B(n26158), .S(gray_img[613]), .O(n26157) );
  MUX2S U30755 ( .A(n15889), .B(n26158), .S(gray_img[608]), .O(n26159) );
  AO12S U30756 ( .B1(n15888), .B2(n26160), .A1(n26159), .O(n14174) );
  INV1S U30757 ( .I(n26169), .O(n26171) );
  MXL2HS U30758 ( .A(gray_img[613]), .B(gray_img[741]), .S(n26198), .OB(n26301) );
  INV1S U30759 ( .I(gray_img[623]), .O(n26183) );
  INV1S U30760 ( .I(gray_img[622]), .O(n26181) );
  INV1S U30761 ( .I(gray_img[621]), .O(n26179) );
  FA1S U30762 ( .A(gray_img[745]), .B(gray_img[744]), .CI(intadd_103_CI), .CO(
        n26175) );
  FA1S U30763 ( .A(n26189), .B(gray_img[746]), .CI(n26175), .CO(n26176) );
  FA1S U30764 ( .A(n26187), .B(gray_img[747]), .CI(n26176), .CO(n26177) );
  FA1S U30765 ( .A(n26185), .B(gray_img[748]), .CI(n26177), .CO(n26178) );
  FA1S U30766 ( .A(n26179), .B(gray_img[749]), .CI(n26178), .CO(n26180) );
  MXL2HS U30767 ( .A(gray_img[621]), .B(gray_img[749]), .S(n26325), .OB(n26195) );
  INV1S U30768 ( .I(gray_img[748]), .O(n26184) );
  MXL2HS U30769 ( .A(n26185), .B(n26184), .S(n26325), .OB(n26303) );
  MXL2HS U30770 ( .A(gray_img[612]), .B(gray_img[740]), .S(n26198), .OB(n26306) );
  INV1S U30771 ( .I(gray_img[747]), .O(n26186) );
  MXL2HS U30772 ( .A(n26187), .B(n26186), .S(n26325), .OB(n26308) );
  MXL2HS U30773 ( .A(gray_img[611]), .B(gray_img[739]), .S(n26198), .OB(n26311) );
  INV1S U30774 ( .I(gray_img[746]), .O(n26188) );
  MXL2HS U30775 ( .A(n26189), .B(n26188), .S(n26325), .OB(n26313) );
  MXL2HS U30776 ( .A(gray_img[610]), .B(gray_img[738]), .S(n26198), .OB(n26316) );
  MXL2HS U30777 ( .A(gray_img[609]), .B(gray_img[737]), .S(n26198), .OB(n26321) );
  MXL2HS U30778 ( .A(gray_img[608]), .B(gray_img[736]), .S(n26198), .OB(n26330) );
  INV1S U30779 ( .I(gray_img[745]), .O(n26190) );
  MXL2HS U30780 ( .A(intadd_103_CI), .B(n26190), .S(n26325), .OB(n26318) );
  INV1S U30781 ( .I(n26196), .O(n26194) );
  NR2 U30782 ( .I1(n26195), .I2(n26194), .O(n26197) );
  INV1S U30783 ( .I(n26195), .O(n26298) );
  OAI22S U30784 ( .A1(n26301), .A2(n26197), .B1(n26196), .B2(n26298), .O(
        n26201) );
  MXL2HS U30785 ( .A(gray_img[622]), .B(gray_img[750]), .S(n26325), .OB(n26208) );
  MXL2HS U30786 ( .A(n26200), .B(n26199), .S(n26198), .OB(n26205) );
  INV1S U30787 ( .I(n26205), .O(n26212) );
  INV1S U30788 ( .I(n26322), .O(n26324) );
  INV1S U30789 ( .I(n26208), .O(n26209) );
  OAI112HS U30790 ( .C1(n26331), .C2(n26212), .A1(n26211), .B1(n26210), .O(
        n14145) );
  MUX2S U30791 ( .A(n15889), .B(n26222), .S(gray_img[869]), .O(n26213) );
  MUX2S U30792 ( .A(n15889), .B(n26222), .S(gray_img[866]), .O(n26216) );
  MUX2S U30793 ( .A(n27447), .B(n26222), .S(gray_img[864]), .O(n26217) );
  AO12S U30794 ( .B1(n15888), .B2(n26224), .A1(n26217), .O(n14130) );
  MUX2S U30795 ( .A(n27447), .B(n27827), .S(gray_img[997]), .O(n26218) );
  MUX2S U30796 ( .A(n27447), .B(n27827), .S(gray_img[994]), .O(n26221) );
  MUX2S U30797 ( .A(n15889), .B(n26222), .S(gray_img[865]), .O(n26223) );
  MUX2S U30798 ( .A(n27447), .B(n27827), .S(gray_img[993]), .O(n26225) );
  INV1S U30799 ( .I(gray_img[877]), .O(n26236) );
  INV1S U30800 ( .I(gray_img[876]), .O(n26232) );
  INV1S U30801 ( .I(gray_img[875]), .O(n26230) );
  INV1S U30802 ( .I(gray_img[874]), .O(n26228) );
  INV1S U30803 ( .I(gray_img[873]), .O(n26226) );
  FA1S U30804 ( .A(gray_img[1001]), .B(gray_img[1000]), .CI(n26226), .CO(
        n26227) );
  FA1S U30805 ( .A(n26228), .B(gray_img[1002]), .CI(n26227), .CO(n26229) );
  FA1S U30806 ( .A(n26230), .B(gray_img[1003]), .CI(n26229), .CO(n26231) );
  INV1S U30807 ( .I(gray_img[1005]), .O(n26233) );
  ND2S U30808 ( .I1(n26233), .I2(gray_img[877]), .O(n26234) );
  AOI22S U30809 ( .A1(gray_img[1005]), .A2(n26236), .B1(n26235), .B2(n26234), 
        .O(n26239) );
  INV1S U30810 ( .I(gray_img[878]), .O(n26237) );
  NR2 U30811 ( .I1(gray_img[1006]), .I2(n26237), .O(n26238) );
  MOAI1S U30812 ( .A1(n26239), .A2(n26238), .B1(gray_img[1006]), .B2(n26237), 
        .O(n26242) );
  ND2S U30813 ( .I1(n26240), .I2(gray_img[879]), .O(n26241) );
  AOI22S U30814 ( .A1(gray_img[1007]), .A2(n26243), .B1(n26242), .B2(n26241), 
        .O(n26256) );
  INV1S U30815 ( .I(gray_img[998]), .O(n26253) );
  INV1S U30816 ( .I(gray_img[997]), .O(n26251) );
  INV1S U30817 ( .I(gray_img[996]), .O(n26249) );
  INV1S U30818 ( .I(gray_img[994]), .O(n26245) );
  FA1S U30819 ( .A(gray_img[865]), .B(gray_img[864]), .CI(intadd_94_CI), .CO(
        n26244) );
  FA1S U30820 ( .A(n26245), .B(gray_img[866]), .CI(n26244), .CO(n26246) );
  FA1S U30821 ( .A(n26247), .B(gray_img[867]), .CI(n26246), .CO(n26248) );
  FA1S U30822 ( .A(n26249), .B(gray_img[868]), .CI(n26248), .CO(n26250) );
  MXL2HS U30823 ( .A(gray_img[998]), .B(gray_img[870]), .S(n27831), .OB(n26269) );
  MXL2HS U30824 ( .A(gray_img[997]), .B(gray_img[869]), .S(n27831), .OB(n26274) );
  MXL2HS U30825 ( .A(gray_img[996]), .B(gray_img[868]), .S(n27831), .OB(n26279) );
  MXL2HS U30826 ( .A(gray_img[995]), .B(gray_img[867]), .S(n27831), .OB(n26284) );
  MXL2HS U30827 ( .A(gray_img[994]), .B(gray_img[866]), .S(n27831), .OB(n26289) );
  MXL2HS U30828 ( .A(gray_img[993]), .B(gray_img[865]), .S(n27831), .OB(n26294) );
  INV1S U30829 ( .I(n26266), .O(n26265) );
  NR2 U30830 ( .I1(n29680), .I2(n26265), .O(n27840) );
  OR2 U30831 ( .I1(n29680), .I2(n26266), .O(n27830) );
  ND2S U30832 ( .I1(n15890), .I2(n27834), .O(n26267) );
  OAI112HS U30833 ( .C1(n27830), .C2(n26269), .A1(n26268), .B1(n26267), .O(
        n26270) );
  OAI112HS U30834 ( .C1(n27830), .C2(n26274), .A1(n26273), .B1(n26272), .O(
        n26275) );
  OAI112HS U30835 ( .C1(n27830), .C2(n26279), .A1(n26278), .B1(n26277), .O(
        n26280) );
  OAI112HS U30836 ( .C1(n27830), .C2(n26284), .A1(n26283), .B1(n26282), .O(
        n26285) );
  OAI112HS U30837 ( .C1(n27830), .C2(n26289), .A1(n26288), .B1(n26287), .O(
        n26290) );
  OAI112HS U30838 ( .C1(n27830), .C2(n26294), .A1(n26293), .B1(n26292), .O(
        n26295) );
  OAI112HS U30839 ( .C1(n26331), .C2(n26301), .A1(n26300), .B1(n26299), .O(
        n14146) );
  OAI112HS U30840 ( .C1(n26331), .C2(n26306), .A1(n26305), .B1(n26304), .O(
        n14147) );
  OAI112HS U30841 ( .C1(n26331), .C2(n26311), .A1(n26310), .B1(n26309), .O(
        n14148) );
  OAI112HS U30842 ( .C1(n26331), .C2(n26316), .A1(n26315), .B1(n26314), .O(
        n14149) );
  OAI112HS U30843 ( .C1(n26331), .C2(n26321), .A1(n26320), .B1(n26319), .O(
        n14150) );
  MUX2S U30844 ( .A(gray_img[616]), .B(gray_img[744]), .S(n26325), .O(n26326)
         );
  OAI112HS U30845 ( .C1(n26331), .C2(n26330), .A1(n26329), .B1(n26328), .O(
        n13780) );
  INV1S U30846 ( .I(gray_img[767]), .O(n26344) );
  INV1S U30847 ( .I(gray_img[764]), .O(n26338) );
  INV1S U30848 ( .I(gray_img[763]), .O(n26336) );
  INV1S U30849 ( .I(gray_img[762]), .O(n26334) );
  MXL2HS U30850 ( .A(gray_img[766]), .B(gray_img[638]), .S(n26480), .OB(n26374) );
  INV1S U30851 ( .I(gray_img[758]), .O(n26354) );
  INV1S U30852 ( .I(gray_img[757]), .O(n26352) );
  INV1S U30853 ( .I(gray_img[756]), .O(n26350) );
  INV1S U30854 ( .I(gray_img[755]), .O(n26348) );
  INV1S U30855 ( .I(gray_img[754]), .O(n26346) );
  FA1S U30856 ( .A(gray_img[625]), .B(gray_img[624]), .CI(intadd_101_CI), .CO(
        n26345) );
  FA1S U30857 ( .A(n26346), .B(gray_img[626]), .CI(n26345), .CO(n26347) );
  FA1S U30858 ( .A(n26348), .B(gray_img[627]), .CI(n26347), .CO(n26349) );
  FA1S U30859 ( .A(n26350), .B(gray_img[628]), .CI(n26349), .CO(n26351) );
  MXL2HS U30860 ( .A(gray_img[765]), .B(gray_img[637]), .S(n26480), .OB(n26448) );
  MXL2HS U30861 ( .A(gray_img[763]), .B(gray_img[635]), .S(n26480), .OB(n26458) );
  MXL2HS U30862 ( .A(gray_img[762]), .B(gray_img[634]), .S(n26480), .OB(n26463) );
  MXL2HS U30863 ( .A(gray_img[761]), .B(gray_img[633]), .S(n26480), .OB(n26476) );
  MXL2HS U30864 ( .A(gray_img[764]), .B(gray_img[636]), .S(n26480), .OB(n26453) );
  NR2 U30865 ( .I1(n26455), .I2(n26453), .O(n26361) );
  OR2 U30866 ( .I1(n29680), .I2(n26368), .O(n26479) );
  INV1S U30867 ( .I(n26368), .O(n26369) );
  OA12S U30868 ( .B1(gray_img[318]), .B2(n29427), .A1(n26483), .O(n26371) );
  MOAI1S U30869 ( .A1(gray_img[318]), .A2(n26483), .B1(n29825), .B2(n26371), 
        .O(n26372) );
  OAI112HS U30870 ( .C1(n26374), .C2(n26479), .A1(n26373), .B1(n26372), .O(
        n14136) );
  FA1S U30871 ( .A(gray_img[1009]), .B(gray_img[1008]), .CI(n26375), .CO(
        n26376) );
  FA1S U30872 ( .A(n26377), .B(gray_img[1010]), .CI(n26376), .CO(n26378) );
  FA1S U30873 ( .A(n26379), .B(gray_img[1011]), .CI(n26378), .CO(n26380) );
  INV1S U30874 ( .I(gray_img[895]), .O(n26400) );
  INV1S U30875 ( .I(gray_img[894]), .O(n26398) );
  INV1S U30876 ( .I(gray_img[893]), .O(n26396) );
  MXL2HS U30877 ( .A(gray_img[894]), .B(gray_img[1022]), .S(n26437), .OB(
        n26414) );
  MXL2HS U30878 ( .A(gray_img[893]), .B(gray_img[1021]), .S(n26437), .OB(
        n26419) );
  MXL2HS U30879 ( .A(gray_img[892]), .B(gray_img[1020]), .S(n26437), .OB(
        n26424) );
  MXL2HS U30880 ( .A(gray_img[891]), .B(gray_img[1019]), .S(n26437), .OB(
        n26429) );
  MXL2HS U30881 ( .A(gray_img[890]), .B(gray_img[1018]), .S(n26437), .OB(
        n26434) );
  MXL2HS U30882 ( .A(gray_img[889]), .B(gray_img[1017]), .S(n26437), .OB(
        n26469) );
  INV1S U30883 ( .I(n26411), .O(n26410) );
  NR2 U30884 ( .I1(n29680), .I2(n26410), .O(n26473) );
  ND2S U30885 ( .I1(n15890), .I2(n26466), .O(n26412) );
  OAI112HS U30886 ( .C1(n26470), .C2(n26414), .A1(n26413), .B1(n26412), .O(
        n26415) );
  OAI112HS U30887 ( .C1(n26470), .C2(n26419), .A1(n26418), .B1(n26417), .O(
        n26420) );
  OAI112HS U30888 ( .C1(n26470), .C2(n26424), .A1(n26423), .B1(n26422), .O(
        n26425) );
  OAI112HS U30889 ( .C1(n26470), .C2(n26429), .A1(n26428), .B1(n26427), .O(
        n26430) );
  OAI112HS U30890 ( .C1(n26470), .C2(n26434), .A1(n26433), .B1(n26432), .O(
        n26435) );
  INV1S U30891 ( .I(n26470), .O(n26439) );
  MUX2S U30892 ( .A(gray_img[888]), .B(gray_img[1016]), .S(n26437), .O(n26438)
         );
  ND2S U30893 ( .I1(n26439), .I2(n26438), .O(n26442) );
  ND2S U30894 ( .I1(n15888), .I2(n26466), .O(n26440) );
  ND3S U30895 ( .I1(n26442), .I2(n26441), .I3(n26440), .O(n26443) );
  ND2S U30896 ( .I1(n26445), .I2(n26483), .O(n26446) );
  OAI112HS U30897 ( .C1(n26479), .C2(n26448), .A1(n26447), .B1(n26446), .O(
        n26449) );
  OAI112HS U30898 ( .C1(n26479), .C2(n26453), .A1(n26452), .B1(n26451), .O(
        n26454) );
  OAI112HS U30899 ( .C1(n26479), .C2(n26458), .A1(n26457), .B1(n26456), .O(
        n26459) );
  OAI112HS U30900 ( .C1(n26479), .C2(n26463), .A1(n26462), .B1(n26461), .O(
        n26464) );
  OAI112HS U30901 ( .C1(n26470), .C2(n26469), .A1(n26468), .B1(n26467), .O(
        n26471) );
  OAI112HS U30902 ( .C1(n26479), .C2(n26476), .A1(n26475), .B1(n26474), .O(
        n26477) );
  INV1S U30903 ( .I(n26479), .O(n26482) );
  MUX2S U30904 ( .A(gray_img[760]), .B(gray_img[632]), .S(n26480), .O(n26481)
         );
  ND2S U30905 ( .I1(n26482), .I2(n26481), .O(n26486) );
  ND2S U30906 ( .I1(n15888), .I2(n26483), .O(n26484) );
  ND3S U30907 ( .I1(n26486), .I2(n26485), .I3(n26484), .O(n26487) );
  INV1S U30908 ( .I(gray_img[318]), .O(n26499) );
  INV1S U30909 ( .I(gray_img[316]), .O(n26495) );
  INV1S U30910 ( .I(gray_img[315]), .O(n26493) );
  INV1S U30911 ( .I(gray_img[314]), .O(n26491) );
  FA1S U30912 ( .A(gray_img[441]), .B(gray_img[440]), .CI(intadd_13_CI), .CO(
        n26490) );
  FA1S U30913 ( .A(n26491), .B(gray_img[442]), .CI(n26490), .CO(n26492) );
  FA1S U30914 ( .A(n26493), .B(gray_img[443]), .CI(n26492), .CO(n26494) );
  FA1S U30915 ( .A(n26495), .B(gray_img[444]), .CI(n26494), .CO(n26496) );
  INV1S U30916 ( .I(gray_img[310]), .O(n26511) );
  INV1S U30917 ( .I(gray_img[309]), .O(n26509) );
  INV1S U30918 ( .I(gray_img[307]), .O(n26505) );
  FA1S U30919 ( .A(intadd_14_CI), .B(gray_img[433]), .CI(intadd_14_B_0_), .CO(
        n26502) );
  MXL2HS U30920 ( .A(gray_img[310]), .B(gray_img[438]), .S(n27842), .OB(n26526) );
  MXL2HS U30921 ( .A(gray_img[309]), .B(gray_img[437]), .S(n27842), .OB(n27796) );
  MXL2HS U30922 ( .A(gray_img[308]), .B(gray_img[436]), .S(n27842), .OB(n27801) );
  MXL2HS U30923 ( .A(gray_img[307]), .B(gray_img[435]), .S(n27842), .OB(n27806) );
  MXL2HS U30924 ( .A(gray_img[306]), .B(gray_img[434]), .S(n27842), .OB(n27811) );
  MXL2HS U30925 ( .A(gray_img[305]), .B(gray_img[433]), .S(n27842), .OB(n27824) );
  INV1S U30926 ( .I(n26523), .O(n26522) );
  NR2 U30927 ( .I1(n29680), .I2(n26522), .O(n27851) );
  OR2 U30928 ( .I1(n29680), .I2(n26523), .O(n27841) );
  ND2S U30929 ( .I1(n15890), .I2(n27845), .O(n26524) );
  OAI112HS U30930 ( .C1(n27841), .C2(n26526), .A1(n26525), .B1(n26524), .O(
        n26527) );
  INV1S U30931 ( .I(gray_img[1567]), .O(n26546) );
  INV1S U30932 ( .I(gray_img[1695]), .O(n26544) );
  INV1S U30933 ( .I(gray_img[1565]), .O(n26529) );
  NR2 U30934 ( .I1(gray_img[1693]), .I2(n26529), .O(n26538) );
  INV1S U30935 ( .I(gray_img[1692]), .O(n26536) );
  INV1S U30936 ( .I(gray_img[1690]), .O(n26532) );
  FA1S U30937 ( .A(gray_img[1561]), .B(gray_img[1560]), .CI(n26530), .CO(
        n26531) );
  FA1S U30938 ( .A(n26532), .B(gray_img[1562]), .CI(n26531), .CO(n26533) );
  FA1S U30939 ( .A(n26534), .B(gray_img[1563]), .CI(n26533), .CO(n26535) );
  MAO222S U30940 ( .A1(gray_img[1564]), .B1(n26536), .C1(n26535), .O(n26537)
         );
  NR2 U30941 ( .I1(n26538), .I2(n26537), .O(n26542) );
  INV1S U30942 ( .I(gray_img[1693]), .O(n26539) );
  INV1S U30943 ( .I(gray_img[1694]), .O(n26540) );
  OAI22S U30944 ( .A1(gray_img[1565]), .A2(n26539), .B1(n26540), .B2(
        gray_img[1566]), .O(n26541) );
  MOAI1S U30945 ( .A1(n26542), .A2(n26541), .B1(gray_img[1566]), .B2(n26540), 
        .O(n26543) );
  OAI12HS U30946 ( .B1(gray_img[1567]), .B2(n26544), .A1(n26543), .O(n26545)
         );
  MXL2HS U30947 ( .A(gray_img[1694]), .B(gray_img[1566]), .S(n26559), .OB(
        n26574) );
  INV1S U30948 ( .I(gray_img[1685]), .O(n26554) );
  INV1S U30949 ( .I(gray_img[1684]), .O(n26552) );
  INV1S U30950 ( .I(gray_img[1683]), .O(n26550) );
  MXL2HS U30951 ( .A(gray_img[1693]), .B(gray_img[1565]), .S(n26559), .OB(
        n29535) );
  MXL2HS U30952 ( .A(gray_img[1692]), .B(gray_img[1564]), .S(n26559), .OB(
        n29540) );
  MUX2S U30953 ( .A(gray_img[1683]), .B(gray_img[1555]), .S(n29577), .O(n29541) );
  MXL2HS U30954 ( .A(gray_img[1691]), .B(gray_img[1563]), .S(n26559), .OB(
        n29545) );
  MUX2S U30955 ( .A(gray_img[1682]), .B(gray_img[1554]), .S(n29577), .O(n29546) );
  MXL2HS U30956 ( .A(gray_img[1690]), .B(gray_img[1562]), .S(n26559), .OB(
        n29550) );
  MXL2HS U30957 ( .A(gray_img[1688]), .B(gray_img[1560]), .S(n26559), .OB(
        n29586) );
  MXL2HS U30958 ( .A(gray_img[1689]), .B(gray_img[1561]), .S(n26559), .OB(
        n29555) );
  MUX2S U30959 ( .A(gray_img[1681]), .B(gray_img[1553]), .S(n29577), .O(n29551) );
  OR2 U30960 ( .I1(n29680), .I2(n26568), .O(n29585) );
  INV1S U30961 ( .I(n26568), .O(n26569) );
  OA12S U30962 ( .B1(gray_img[782]), .B2(n29427), .A1(n29580), .O(n26571) );
  MOAI1S U30963 ( .A1(gray_img[782]), .A2(n29580), .B1(n29825), .B2(n26571), 
        .O(n26572) );
  OAI112HS U30964 ( .C1(n26574), .C2(n29585), .A1(n26573), .B1(n26572), .O(
        n13897) );
  INV1S U30965 ( .I(gray_img[1678]), .O(n26585) );
  INV1S U30966 ( .I(gray_img[1677]), .O(n26583) );
  INV1S U30967 ( .I(gray_img[1675]), .O(n26579) );
  FA1S U30968 ( .A(gray_img[1545]), .B(gray_img[1544]), .CI(n26575), .CO(
        n26576) );
  FA1S U30969 ( .A(n26590), .B(gray_img[1666]), .CI(n26589), .CO(n26591) );
  FA1S U30970 ( .A(n26592), .B(gray_img[1667]), .CI(n26591), .CO(n26593) );
  MXL2HS U30971 ( .A(gray_img[1542]), .B(gray_img[1670]), .S(n29478), .OB(
        n26614) );
  MXL2HS U30972 ( .A(gray_img[1541]), .B(gray_img[1669]), .S(n29478), .OB(
        n29434) );
  MXL2HS U30973 ( .A(gray_img[1540]), .B(gray_img[1668]), .S(n29478), .OB(
        n29439) );
  MXL2HS U30974 ( .A(gray_img[1539]), .B(gray_img[1667]), .S(n29478), .OB(
        n29444) );
  MUX2S U30975 ( .A(gray_img[1674]), .B(gray_img[1546]), .S(n26601), .O(n29451) );
  MXL2HS U30976 ( .A(gray_img[1538]), .B(gray_img[1666]), .S(n29478), .OB(
        n29449) );
  MUX2S U30977 ( .A(gray_img[1673]), .B(gray_img[1545]), .S(n26601), .O(n29456) );
  MXL2HS U30978 ( .A(gray_img[1537]), .B(gray_img[1665]), .S(n29478), .OB(
        n29454) );
  MUX2S U30979 ( .A(gray_img[1672]), .B(gray_img[1544]), .S(n26601), .O(n29486) );
  INV1S U30980 ( .I(n26611), .O(n26610) );
  NR2 U30981 ( .I1(n29680), .I2(n26610), .O(n29487) );
  ND2S U30982 ( .I1(n15890), .I2(n29481), .O(n26612) );
  OAI112HS U30983 ( .C1(n29477), .C2(n26614), .A1(n26613), .B1(n26612), .O(
        n26615) );
  MAO222S U30984 ( .A1(gray_img[1161]), .B1(gray_img[1160]), .C1(intadd_89_CI), 
        .O(n26617) );
  FA1S U30985 ( .A(intadd_89_B_1_), .B(gray_img[1162]), .CI(n26617), .CO(
        n26618) );
  FA1S U30986 ( .A(n26619), .B(gray_img[1163]), .CI(n26618), .CO(n26620) );
  MXL2HS U30987 ( .A(gray_img[1038]), .B(gray_img[1166]), .S(n26640), .OB(
        n26655) );
  INV1S U30988 ( .I(gray_img[1157]), .O(n26635) );
  MAO222S U30989 ( .A1(gray_img[1025]), .B1(gray_img[1024]), .C1(intadd_88_CI), 
        .O(n26628) );
  FA1S U30990 ( .A(n26629), .B(gray_img[1026]), .CI(n26628), .CO(n26630) );
  FA1S U30991 ( .A(n26631), .B(gray_img[1027]), .CI(n26630), .CO(n26632) );
  FA1S U30992 ( .A(n26633), .B(gray_img[1028]), .CI(n26632), .CO(n26634) );
  MXL2HS U30993 ( .A(gray_img[1037]), .B(gray_img[1165]), .S(n26640), .OB(
        n29715) );
  MXL2HS U30994 ( .A(gray_img[1036]), .B(gray_img[1164]), .S(n26640), .OB(
        n29720) );
  MXL2HS U30995 ( .A(gray_img[1035]), .B(gray_img[1163]), .S(n26640), .OB(
        n29725) );
  MXL2HS U30996 ( .A(gray_img[1034]), .B(gray_img[1162]), .S(n26640), .OB(
        n29730) );
  MXL2HS U30997 ( .A(gray_img[1032]), .B(gray_img[1160]), .S(n26640), .OB(
        n29737) );
  MXL2HS U30998 ( .A(gray_img[1033]), .B(gray_img[1161]), .S(n26640), .OB(
        n29746) );
  MUX2S U30999 ( .A(gray_img[1153]), .B(gray_img[1025]), .S(n29731), .O(n29738) );
  OR2 U31000 ( .I1(n29680), .I2(n26649), .O(n29745) );
  INV1S U31001 ( .I(n26649), .O(n26650) );
  OA12S U31002 ( .B1(gray_img[518]), .B2(n29427), .A1(n29740), .O(n26652) );
  MOAI1S U31003 ( .A1(gray_img[518]), .A2(n29740), .B1(n29825), .B2(n26652), 
        .O(n26653) );
  OAI112HS U31004 ( .C1(n26655), .C2(n29745), .A1(n26654), .B1(n26653), .O(
        n14067) );
  FA1S U31005 ( .A(n26656), .B(intadd_28_A_0_), .CI(gray_img[1825]), .CO(
        n26657) );
  FA1S U31006 ( .A(gray_img[1826]), .B(n26658), .CI(n26657), .CO(n26659) );
  FA1S U31007 ( .A(gray_img[1827]), .B(n26660), .CI(n26659), .CO(n26661) );
  MXL2HS U31008 ( .A(gray_img[1958]), .B(gray_img[1830]), .S(n26682), .OB(
        n26697) );
  FA1S U31009 ( .A(gray_img[1833]), .B(gray_img[1832]), .CI(n26669), .CO(
        n26670) );
  FA1S U31010 ( .A(n26671), .B(gray_img[1834]), .CI(n26670), .CO(n26672) );
  FA1S U31011 ( .A(n26673), .B(gray_img[1835]), .CI(n26672), .CO(n26674) );
  MXL2HS U31012 ( .A(gray_img[1957]), .B(gray_img[1829]), .S(n26682), .OB(
        n29166) );
  MXL2HS U31013 ( .A(gray_img[1956]), .B(gray_img[1828]), .S(n26682), .OB(
        n29171) );
  MXL2HS U31014 ( .A(gray_img[1955]), .B(gray_img[1827]), .S(n26682), .OB(
        n29176) );
  MXL2HS U31015 ( .A(gray_img[1954]), .B(gray_img[1826]), .S(n26682), .OB(
        n29181) );
  MXL2HS U31016 ( .A(gray_img[1953]), .B(gray_img[1825]), .S(n26682), .OB(
        n29197) );
  MXL2HS U31017 ( .A(gray_img[1952]), .B(gray_img[1824]), .S(n26682), .OB(
        n30027) );
  OR2 U31018 ( .I1(n29680), .I2(n26691), .O(n30026) );
  INV1S U31019 ( .I(n26691), .O(n26692) );
  OA12S U31020 ( .B1(gray_img[918]), .B2(n29427), .A1(n30021), .O(n26694) );
  MOAI1S U31021 ( .A1(n30021), .A2(gray_img[918]), .B1(n29825), .B2(n26694), 
        .O(n26695) );
  OAI112HS U31022 ( .C1(n26697), .C2(n30026), .A1(n26696), .B1(n26695), .O(
        n13829) );
  MUX2S U31023 ( .A(n27447), .B(n26707), .S(gray_img[92]), .O(n26699) );
  MUX2S U31024 ( .A(n27447), .B(n26707), .S(gray_img[90]), .O(n26701) );
  MUX2S U31025 ( .A(n27447), .B(n26707), .S(gray_img[88]), .O(n26702) );
  AO12S U31026 ( .B1(n19092), .B2(n26709), .A1(n26702), .O(n14263) );
  MUX2S U31027 ( .A(n27447), .B(n26724), .S(gray_img[221]), .O(n26703) );
  MUX2S U31028 ( .A(n27447), .B(n26724), .S(gray_img[218]), .O(n26706) );
  MUX2S U31029 ( .A(n28534), .B(n26724), .S(gray_img[217]), .O(n26710) );
  AO12S U31030 ( .B1(n15891), .B2(n26722), .A1(n26711), .O(n15266) );
  MUX2S U31031 ( .A(n27447), .B(n26720), .S(gray_img[84]), .O(n26712) );
  MUX2S U31032 ( .A(n27447), .B(n26720), .S(gray_img[82]), .O(n26714) );
  MUX2S U31033 ( .A(n27447), .B(n26839), .S(gray_img[213]), .O(n26716) );
  MUX2S U31034 ( .A(n27447), .B(n26839), .S(gray_img[212]), .O(n26717) );
  MUX2S U31035 ( .A(n27447), .B(n26839), .S(gray_img[211]), .O(n26718) );
  MUX2S U31036 ( .A(n27447), .B(n26839), .S(gray_img[210]), .O(n26719) );
  MUX2S U31037 ( .A(n27447), .B(n26839), .S(gray_img[209]), .O(n26723) );
  MUX2S U31038 ( .A(n15889), .B(n26724), .S(gray_img[216]), .O(n26725) );
  AO12S U31039 ( .B1(n15888), .B2(n26726), .A1(n26725), .O(n14248) );
  ND2S U31040 ( .I1(n15890), .I2(n26842), .O(n26727) );
  OAI112HS U31041 ( .C1(n26846), .C2(n26729), .A1(n26728), .B1(n26727), .O(
        n26730) );
  MUX2S U31042 ( .A(n27447), .B(n26741), .S(gray_img[340]), .O(n26733) );
  MUX2S U31043 ( .A(n27447), .B(n26745), .S(gray_img[465]), .O(n26740) );
  AO12S U31044 ( .B1(n19092), .B2(n26743), .A1(n26742), .O(n14220) );
  MUX2S U31045 ( .A(n27447), .B(n26745), .S(gray_img[464]), .O(n26746) );
  AO12S U31046 ( .B1(n15888), .B2(n26747), .A1(n26746), .O(n14205) );
  MUX2S U31047 ( .A(n27447), .B(n26757), .S(gray_img[349]), .O(n26748) );
  MUX2S U31048 ( .A(n27447), .B(n26757), .S(gray_img[347]), .O(n26750) );
  MUX2S U31049 ( .A(n28534), .B(n26757), .S(gray_img[346]), .O(n26751) );
  AO12S U31050 ( .B1(n19092), .B2(n26759), .A1(n26752), .O(n14219) );
  MUX2S U31051 ( .A(n27447), .B(n27350), .S(gray_img[476]), .O(n26754) );
  MUX2S U31052 ( .A(n27447), .B(n27350), .S(gray_img[475]), .O(n26755) );
  MUX2S U31053 ( .A(n28534), .B(n27350), .S(gray_img[474]), .O(n26756) );
  INV1S U31054 ( .I(gray_img[343]), .O(n26774) );
  INV1S U31055 ( .I(gray_img[342]), .O(n26772) );
  INV1S U31056 ( .I(gray_img[341]), .O(n26770) );
  INV1S U31057 ( .I(gray_img[340]), .O(n26768) );
  INV1S U31058 ( .I(gray_img[339]), .O(n26766) );
  INV1S U31059 ( .I(gray_img[337]), .O(n26761) );
  NR2 U31060 ( .I1(gray_img[465]), .I2(n26761), .O(n26762) );
  MOAI1S U31061 ( .A1(n26762), .A2(gray_img[336]), .B1(n26761), .B2(
        gray_img[465]), .O(n26764) );
  INV1S U31062 ( .I(gray_img[338]), .O(n26763) );
  MXL2HS U31063 ( .A(gray_img[342]), .B(gray_img[470]), .S(n26787), .OB(n26802) );
  INV1S U31064 ( .I(gray_img[478]), .O(n26784) );
  INV1S U31065 ( .I(gray_img[477]), .O(n26782) );
  INV1S U31066 ( .I(gray_img[476]), .O(n26780) );
  INV1S U31067 ( .I(gray_img[475]), .O(n26778) );
  INV1S U31068 ( .I(gray_img[474]), .O(n26776) );
  MAO222S U31069 ( .A1(gray_img[345]), .B1(gray_img[344]), .C1(intadd_117_CI), 
        .O(n26775) );
  FA1S U31070 ( .A(n26776), .B(gray_img[346]), .CI(n26775), .CO(n26777) );
  FA1S U31071 ( .A(n26778), .B(gray_img[347]), .CI(n26777), .CO(n26779) );
  FA1S U31072 ( .A(n26780), .B(gray_img[348]), .CI(n26779), .CO(n26781) );
  MAO222 U31073 ( .A1(n26786), .B1(gray_img[351]), .C1(n26785), .O(n27353) );
  MXL2HS U31074 ( .A(gray_img[341]), .B(gray_img[469]), .S(n26787), .OB(n26807) );
  MXL2HS U31075 ( .A(gray_img[340]), .B(gray_img[468]), .S(n26787), .OB(n26812) );
  MXL2HS U31076 ( .A(gray_img[339]), .B(gray_img[467]), .S(n26787), .OB(n26817) );
  MXL2HS U31077 ( .A(gray_img[338]), .B(gray_img[466]), .S(n26787), .OB(n26822) );
  MXL2HS U31078 ( .A(gray_img[337]), .B(gray_img[465]), .S(n26787), .OB(n26827) );
  MXL2HS U31079 ( .A(gray_img[336]), .B(gray_img[464]), .S(n26787), .OB(n27362) );
  OR2 U31080 ( .I1(n29680), .I2(n26796), .O(n27361) );
  INV1S U31081 ( .I(n26796), .O(n26797) );
  ND2S U31082 ( .I1(n27355), .I2(n26798), .O(n26801) );
  INV1S U31083 ( .I(n27356), .O(n27358) );
  OAI112HS U31084 ( .C1(n26802), .C2(n27361), .A1(n26801), .B1(n26800), .O(
        n14198) );
  ND2S U31085 ( .I1(n27355), .I2(n26803), .O(n26806) );
  MUX2S U31086 ( .A(n30005), .B(n27356), .S(gray_img[173]), .O(n26804) );
  OA12S U31087 ( .B1(n29831), .B2(n27358), .A1(n26804), .O(n26805) );
  OAI112HS U31088 ( .C1(n26807), .C2(n27361), .A1(n26806), .B1(n26805), .O(
        n14199) );
  ND2S U31089 ( .I1(n27355), .I2(n26808), .O(n26811) );
  OAI112HS U31090 ( .C1(n26812), .C2(n27361), .A1(n26811), .B1(n26810), .O(
        n14200) );
  ND2S U31091 ( .I1(n27355), .I2(n26813), .O(n26816) );
  OAI112HS U31092 ( .C1(n26817), .C2(n27361), .A1(n26816), .B1(n26815), .O(
        n14201) );
  ND2S U31093 ( .I1(n27355), .I2(n26818), .O(n26821) );
  OAI112HS U31094 ( .C1(n26822), .C2(n27361), .A1(n26821), .B1(n26820), .O(
        n14202) );
  ND2S U31095 ( .I1(n27355), .I2(n26823), .O(n26826) );
  MUX2S U31096 ( .A(n30005), .B(n27356), .S(gray_img[169]), .O(n26824) );
  OA12S U31097 ( .B1(n29884), .B2(n27358), .A1(n26824), .O(n26825) );
  OAI112HS U31098 ( .C1(n26827), .C2(n27361), .A1(n26826), .B1(n26825), .O(
        n14203) );
  ND2S U31099 ( .I1(n26828), .I2(n26842), .O(n26829) );
  OAI112HS U31100 ( .C1(n26846), .C2(n26831), .A1(n26830), .B1(n26829), .O(
        n26832) );
  OAI112HS U31101 ( .C1(n26846), .C2(n26836), .A1(n26835), .B1(n26834), .O(
        n26837) );
  MUX2S U31102 ( .A(n27447), .B(n26839), .S(gray_img[208]), .O(n26840) );
  AO12S U31103 ( .B1(n15888), .B2(n26841), .A1(n26840), .O(n14249) );
  ND2S U31104 ( .I1(n15928), .I2(n26842), .O(n26843) );
  OAI112HS U31105 ( .C1(n26846), .C2(n26845), .A1(n26844), .B1(n26843), .O(
        n26847) );
  MUX2S U31106 ( .A(n15889), .B(n26859), .S(gray_img[333]), .O(n26850) );
  MUX2S U31107 ( .A(n15889), .B(n26859), .S(gray_img[332]), .O(n26851) );
  MUX2S U31108 ( .A(n15889), .B(n26859), .S(gray_img[331]), .O(n26852) );
  MUX2S U31109 ( .A(n15889), .B(n26859), .S(gray_img[330]), .O(n26853) );
  MUX2S U31110 ( .A(n15889), .B(n26859), .S(gray_img[328]), .O(n26854) );
  AO12S U31111 ( .B1(n15888), .B2(n26861), .A1(n26854), .O(n14221) );
  MUX2S U31112 ( .A(n15889), .B(n26940), .S(gray_img[460]), .O(n26856) );
  MUX2S U31113 ( .A(n15889), .B(n26940), .S(gray_img[459]), .O(n26857) );
  MUX2S U31114 ( .A(n15889), .B(n26940), .S(gray_img[458]), .O(n26858) );
  ND2S U31115 ( .I1(n15890), .I2(n26932), .O(n26863) );
  OAI112HS U31116 ( .C1(n26936), .C2(n26865), .A1(n26864), .B1(n26863), .O(
        n26866) );
  MUX2S U31117 ( .A(n27447), .B(n26877), .S(gray_img[76]), .O(n26869) );
  MUX2S U31118 ( .A(n28534), .B(n26877), .S(gray_img[74]), .O(n26871) );
  AO12S U31119 ( .B1(n15888), .B2(n26879), .A1(n26872), .O(n14265) );
  MUX2S U31120 ( .A(n15889), .B(n26881), .S(gray_img[205]), .O(n26873) );
  MUX2S U31121 ( .A(n27447), .B(n26881), .S(gray_img[204]), .O(n26874) );
  MUX2S U31122 ( .A(n15889), .B(n26881), .S(gray_img[202]), .O(n26876) );
  MUX2S U31123 ( .A(n15889), .B(n26881), .S(gray_img[201]), .O(n26880) );
  MUX2S U31124 ( .A(n15889), .B(n26881), .S(gray_img[200]), .O(n26882) );
  AO12S U31125 ( .B1(n15888), .B2(n26883), .A1(n26882), .O(n14257) );
  OAI112HS U31126 ( .C1(n26928), .C2(n26886), .A1(n26885), .B1(n26884), .O(
        n26887) );
  OAI112HS U31127 ( .C1(n26928), .C2(n26891), .A1(n26890), .B1(n26889), .O(
        n26892) );
  OAI112HS U31128 ( .C1(n26928), .C2(n26896), .A1(n26895), .B1(n26894), .O(
        n26897) );
  OAI112HS U31129 ( .C1(n26928), .C2(n26901), .A1(n26900), .B1(n26899), .O(
        n26902) );
  OAI112HS U31130 ( .C1(n26936), .C2(n26906), .A1(n26905), .B1(n26904), .O(
        n26907) );
  OAI112HS U31131 ( .C1(n26936), .C2(n26911), .A1(n26910), .B1(n26909), .O(
        n26912) );
  OAI112HS U31132 ( .C1(n26936), .C2(n26916), .A1(n26915), .B1(n26914), .O(
        n26917) );
  OAI112HS U31133 ( .C1(n26936), .C2(n26921), .A1(n26920), .B1(n26919), .O(
        n26922) );
  OAI112HS U31134 ( .C1(n26928), .C2(n26927), .A1(n26926), .B1(n26925), .O(
        n26929) );
  OAI112HS U31135 ( .C1(n26936), .C2(n26935), .A1(n26934), .B1(n26933), .O(
        n26937) );
  AO12S U31136 ( .B1(n15888), .B2(n26942), .A1(n26941), .O(n14213) );
  INV1S U31137 ( .I(gray_img[166]), .O(n26953) );
  INV1S U31138 ( .I(gray_img[165]), .O(n26951) );
  INV1S U31139 ( .I(gray_img[164]), .O(n26949) );
  INV1S U31140 ( .I(gray_img[163]), .O(n26947) );
  INV1S U31141 ( .I(gray_img[162]), .O(n26945) );
  INV1S U31142 ( .I(gray_img[161]), .O(n26943) );
  FA1S U31143 ( .A(n26945), .B(gray_img[34]), .CI(n26944), .CO(n26946) );
  INV1S U31144 ( .I(gray_img[45]), .O(n26964) );
  INV1S U31145 ( .I(gray_img[44]), .O(n26962) );
  MXL2HS U31146 ( .A(gray_img[46]), .B(gray_img[174]), .S(n27363), .OB(n26982)
         );
  MXL2HS U31147 ( .A(gray_img[45]), .B(gray_img[173]), .S(n27363), .OB(n27332)
         );
  MXL2HS U31148 ( .A(gray_img[44]), .B(gray_img[172]), .S(n27363), .OB(n27337)
         );
  MXL2HS U31149 ( .A(gray_img[43]), .B(gray_img[171]), .S(n27363), .OB(n27342)
         );
  MXL2HS U31150 ( .A(gray_img[42]), .B(gray_img[170]), .S(n27363), .OB(n27347)
         );
  MUX2S U31151 ( .A(gray_img[160]), .B(gray_img[32]), .S(n26969), .O(n27370)
         );
  MXL2HS U31152 ( .A(gray_img[41]), .B(gray_img[169]), .S(n27363), .OB(n27374)
         );
  INV1S U31153 ( .I(n26979), .O(n26978) );
  NR2 U31154 ( .I1(n29680), .I2(n26978), .O(n27378) );
  OR2 U31155 ( .I1(n29680), .I2(n26979), .O(n27375) );
  ND2S U31156 ( .I1(n15890), .I2(n27371), .O(n26980) );
  OAI112HS U31157 ( .C1(n27375), .C2(n26982), .A1(n26981), .B1(n26980), .O(
        n26983) );
  MUX2S U31158 ( .A(n15889), .B(n26994), .S(gray_img[732]), .O(n26986) );
  MUX2S U31159 ( .A(n15889), .B(n26994), .S(gray_img[731]), .O(n26987) );
  MUX2S U31160 ( .A(n15889), .B(n26994), .S(gray_img[728]), .O(n26989) );
  AO12S U31161 ( .B1(n15888), .B2(n26996), .A1(n26989), .O(n14160) );
  MUX2S U31162 ( .A(n27447), .B(n27103), .S(gray_img[605]), .O(n26990) );
  MUX2S U31163 ( .A(n27447), .B(n27103), .S(gray_img[604]), .O(n26991) );
  MUX2S U31164 ( .A(n27447), .B(n26994), .S(gray_img[729]), .O(n26995) );
  MUX2S U31165 ( .A(n27447), .B(n27007), .S(gray_img[725]), .O(n26998) );
  MUX2S U31166 ( .A(n15889), .B(n27007), .S(gray_img[723]), .O(n27000) );
  MUX2S U31167 ( .A(n15889), .B(n27007), .S(gray_img[722]), .O(n27001) );
  MUX2S U31168 ( .A(n15889), .B(n27007), .S(gray_img[720]), .O(n27002) );
  AO12S U31169 ( .B1(n19092), .B2(n27009), .A1(n27002), .O(n14161) );
  MUX2S U31170 ( .A(n27447), .B(n27011), .S(gray_img[597]), .O(n27003) );
  MUX2S U31171 ( .A(n15889), .B(n27011), .S(gray_img[592]), .O(n27012) );
  AO12S U31172 ( .B1(n15888), .B2(n27013), .A1(n27012), .O(n14176) );
  INV1S U31173 ( .I(gray_img[607]), .O(n27037) );
  INV1S U31174 ( .I(gray_img[606]), .O(n27035) );
  INV1S U31175 ( .I(gray_img[602]), .O(n27027) );
  FA1S U31176 ( .A(gray_img[729]), .B(gray_img[728]), .CI(intadd_106_CI), .CO(
        n27026) );
  FA1S U31177 ( .A(n27027), .B(gray_img[730]), .CI(n27026), .CO(n27028) );
  FA1S U31178 ( .A(n27029), .B(gray_img[731]), .CI(n27028), .CO(n27030) );
  FA1S U31179 ( .A(n27031), .B(gray_img[732]), .CI(n27030), .CO(n27032) );
  FA1S U31180 ( .A(n27033), .B(gray_img[733]), .CI(n27032), .CO(n27034) );
  MXL2HS U31181 ( .A(gray_img[606]), .B(gray_img[734]), .S(n27106), .OB(n27051) );
  MXL2HS U31182 ( .A(gray_img[605]), .B(gray_img[733]), .S(n27106), .OB(n27085) );
  MXL2HS U31183 ( .A(gray_img[604]), .B(gray_img[732]), .S(n27106), .OB(n27090) );
  MXL2HS U31184 ( .A(gray_img[603]), .B(gray_img[731]), .S(n27106), .OB(n27095) );
  MXL2HS U31185 ( .A(gray_img[602]), .B(gray_img[730]), .S(n27106), .OB(n27100) );
  MXL2HS U31186 ( .A(gray_img[601]), .B(gray_img[729]), .S(n27106), .OB(n27117) );
  MAO222 U31187 ( .A1(n27113), .B1(n27117), .C1(n27120), .O(n27039) );
  MAO222 U31188 ( .A1(n27046), .B1(n27045), .C1(n27044), .O(n27048) );
  INV1S U31189 ( .I(n27048), .O(n27047) );
  NR2 U31190 ( .I1(n29680), .I2(n27047), .O(n27121) );
  OR2 U31191 ( .I1(n29680), .I2(n27048), .O(n27118) );
  ND2S U31192 ( .I1(n15890), .I2(n27114), .O(n27049) );
  OAI112HS U31193 ( .C1(n27118), .C2(n27051), .A1(n27050), .B1(n27049), .O(
        n27052) );
  MUX2S U31194 ( .A(n15889), .B(n27063), .S(gray_img[981]), .O(n27054) );
  MUX2S U31195 ( .A(n27447), .B(n27063), .S(gray_img[979]), .O(n27056) );
  MUX2S U31196 ( .A(n15889), .B(n27063), .S(gray_img[978]), .O(n27057) );
  MUX2S U31197 ( .A(n15889), .B(n27063), .S(gray_img[976]), .O(n27058) );
  AO12S U31198 ( .B1(n15888), .B2(n27065), .A1(n27058), .O(n14117) );
  MUX2S U31199 ( .A(n15889), .B(n27067), .S(gray_img[853]), .O(n27059) );
  MUX2S U31200 ( .A(n15889), .B(n27067), .S(gray_img[852]), .O(n27060) );
  MUX2S U31201 ( .A(n27447), .B(n27067), .S(gray_img[851]), .O(n27061) );
  MUX2S U31202 ( .A(n15889), .B(n27067), .S(gray_img[850]), .O(n27062) );
  MUX2S U31203 ( .A(n15889), .B(n27063), .S(gray_img[977]), .O(n27064) );
  MUX2S U31204 ( .A(n15889), .B(n27067), .S(gray_img[849]), .O(n27066) );
  MUX2S U31205 ( .A(n27447), .B(n27067), .S(gray_img[848]), .O(n27068) );
  AO12S U31206 ( .B1(n15888), .B2(n27069), .A1(n27068), .O(n14132) );
  MUX2S U31207 ( .A(n27447), .B(n27079), .S(gray_img[989]), .O(n27070) );
  MUX2S U31208 ( .A(n15889), .B(n27079), .S(gray_img[988]), .O(n27071) );
  MUX2S U31209 ( .A(n15889), .B(n27079), .S(gray_img[987]), .O(n27072) );
  MUX2S U31210 ( .A(n15889), .B(n27079), .S(gray_img[986]), .O(n27073) );
  MUX2S U31211 ( .A(n15889), .B(n27079), .S(gray_img[984]), .O(n27074) );
  AO12S U31212 ( .B1(n19092), .B2(n27081), .A1(n27074), .O(n14116) );
  MUX2S U31213 ( .A(n15889), .B(n30063), .S(gray_img[860]), .O(n27076) );
  MUX2S U31214 ( .A(n15889), .B(n30063), .S(gray_img[859]), .O(n27077) );
  MUX2S U31215 ( .A(n15889), .B(n30063), .S(gray_img[858]), .O(n27078) );
  MUX2S U31216 ( .A(n27447), .B(n27079), .S(gray_img[985]), .O(n27080) );
  MUX2S U31217 ( .A(n15889), .B(n30063), .S(gray_img[857]), .O(n27082) );
  OAI112HS U31218 ( .C1(n27118), .C2(n27085), .A1(n27084), .B1(n27083), .O(
        n27086) );
  OAI112HS U31219 ( .C1(n27118), .C2(n27090), .A1(n27089), .B1(n27088), .O(
        n27091) );
  OAI112HS U31220 ( .C1(n27118), .C2(n27095), .A1(n27094), .B1(n27093), .O(
        n27096) );
  OAI112HS U31221 ( .C1(n27118), .C2(n27100), .A1(n27099), .B1(n27098), .O(
        n27101) );
  AO12S U31222 ( .B1(n15888), .B2(n27105), .A1(n27104), .O(n14175) );
  INV1S U31223 ( .I(n27118), .O(n27108) );
  MUX2S U31224 ( .A(gray_img[600]), .B(gray_img[728]), .S(n27106), .O(n27107)
         );
  ND2S U31225 ( .I1(n27108), .I2(n27107), .O(n27111) );
  ND2S U31226 ( .I1(n15888), .I2(n27114), .O(n27109) );
  ND3S U31227 ( .I1(n27111), .I2(n27110), .I3(n27109), .O(n27112) );
  OAI112HS U31228 ( .C1(n27118), .C2(n27117), .A1(n27116), .B1(n27115), .O(
        n27119) );
  MUX2S U31229 ( .A(n15889), .B(n27131), .S(gray_img[587]), .O(n27124) );
  MUX2S U31230 ( .A(n15889), .B(n27131), .S(gray_img[586]), .O(n27125) );
  MUX2S U31231 ( .A(n15889), .B(n27131), .S(gray_img[584]), .O(n27126) );
  AO12S U31232 ( .B1(n15888), .B2(n27133), .A1(n27126), .O(n14177) );
  MUX2S U31233 ( .A(n15889), .B(n27241), .S(gray_img[716]), .O(n27128) );
  MUX2S U31234 ( .A(n15889), .B(n27241), .S(gray_img[715]), .O(n27129) );
  MUX2S U31235 ( .A(n15889), .B(n27241), .S(gray_img[714]), .O(n27130) );
  MUX2S U31236 ( .A(n15889), .B(n27131), .S(gray_img[585]), .O(n27132) );
  MUX2S U31237 ( .A(n27447), .B(n27241), .S(gray_img[713]), .O(n27134) );
  FA1S U31238 ( .A(gray_img[577]), .B(gray_img[576]), .CI(intadd_109_CI), .CO(
        n27135) );
  FA1S U31239 ( .A(n27136), .B(gray_img[578]), .CI(n27135), .CO(n27137) );
  FA1S U31240 ( .A(n27138), .B(gray_img[579]), .CI(n27137), .CO(n27139) );
  MXL2HS U31241 ( .A(gray_img[710]), .B(gray_img[582]), .S(n27159), .OB(n27174) );
  INV1S U31242 ( .I(gray_img[718]), .O(n27156) );
  INV1S U31243 ( .I(gray_img[717]), .O(n27154) );
  INV1S U31244 ( .I(gray_img[716]), .O(n27152) );
  INV1S U31245 ( .I(gray_img[715]), .O(n27150) );
  INV1S U31246 ( .I(gray_img[714]), .O(n27148) );
  FA1S U31247 ( .A(gray_img[585]), .B(gray_img[584]), .CI(intadd_108_CI), .CO(
        n27147) );
  FA1S U31248 ( .A(n27148), .B(gray_img[586]), .CI(n27147), .CO(n27149) );
  MXL2HS U31249 ( .A(gray_img[709]), .B(gray_img[581]), .S(n27159), .OB(n27206) );
  MXL2HS U31250 ( .A(gray_img[708]), .B(gray_img[580]), .S(n27159), .OB(n27211) );
  MXL2HS U31251 ( .A(gray_img[707]), .B(gray_img[579]), .S(n27159), .OB(n27235) );
  MXL2HS U31252 ( .A(gray_img[706]), .B(gray_img[578]), .S(n27159), .OB(n27240) );
  MXL2HS U31253 ( .A(gray_img[705]), .B(gray_img[577]), .S(n27159), .OB(n27258) );
  MXL2HS U31254 ( .A(gray_img[704]), .B(gray_img[576]), .S(n27159), .OB(n27249) );
  OR2 U31255 ( .I1(n29680), .I2(n27168), .O(n27257) );
  INV1S U31256 ( .I(n27168), .O(n27169) );
  OAI112HS U31257 ( .C1(n27174), .C2(n27257), .A1(n27173), .B1(n27172), .O(
        n14163) );
  ND2S U31258 ( .I1(n27259), .I2(gray_img[973]), .O(n27177) );
  ND2S U31259 ( .I1(n27447), .I2(n27175), .O(n27176) );
  OAI112HS U31260 ( .C1(n29831), .C2(n27259), .A1(n27177), .B1(n27176), .O(
        n15211) );
  ND2S U31261 ( .I1(n27188), .I2(gray_img[845]), .O(n27180) );
  ND2S U31262 ( .I1(n27447), .I2(n27178), .O(n27179) );
  OAI112HS U31263 ( .C1(n29831), .C2(n27188), .A1(n27180), .B1(n27179), .O(
        n15219) );
  MUX2S U31264 ( .A(n15889), .B(n27188), .S(gray_img[843]), .O(n27182) );
  MUX2S U31265 ( .A(n15889), .B(n27188), .S(gray_img[842]), .O(n27183) );
  MUX2S U31266 ( .A(n15889), .B(n27188), .S(gray_img[840]), .O(n27184) );
  AO12S U31267 ( .B1(n15888), .B2(n27190), .A1(n27184), .O(n14133) );
  MUX2S U31268 ( .A(n15889), .B(n27259), .S(gray_img[971]), .O(n27186) );
  MUX2S U31269 ( .A(n15889), .B(n27259), .S(gray_img[970]), .O(n27187) );
  MUX2S U31270 ( .A(n15889), .B(n27188), .S(gray_img[841]), .O(n27189) );
  OAI112HS U31271 ( .C1(n27230), .C2(n27196), .A1(n27195), .B1(n27194), .O(
        n14119) );
  OAI112HS U31272 ( .C1(n27230), .C2(n27201), .A1(n27200), .B1(n27199), .O(
        n14121) );
  OAI112HS U31273 ( .C1(n27206), .C2(n27257), .A1(n27205), .B1(n27204), .O(
        n14164) );
  OAI112HS U31274 ( .C1(n27211), .C2(n27257), .A1(n27210), .B1(n27209), .O(
        n14165) );
  OAI112HS U31275 ( .C1(n27230), .C2(n27216), .A1(n27215), .B1(n27214), .O(
        n14122) );
  OAI112HS U31276 ( .C1(n27230), .C2(n27221), .A1(n27220), .B1(n27219), .O(
        n14123) );
  OAI112HS U31277 ( .C1(n27230), .C2(n27229), .A1(n27228), .B1(n27227), .O(
        n14124) );
  OAI112HS U31278 ( .C1(n27235), .C2(n27257), .A1(n27234), .B1(n27233), .O(
        n14166) );
  OAI112HS U31279 ( .C1(n27240), .C2(n27257), .A1(n27239), .B1(n27238), .O(
        n14167) );
  MUX2S U31280 ( .A(n15889), .B(n27241), .S(gray_img[712]), .O(n27242) );
  AO12S U31281 ( .B1(n15888), .B2(n27243), .A1(n27242), .O(n14169) );
  MUX2S U31282 ( .A(gray_img[712]), .B(gray_img[584]), .S(n27244), .O(n27245)
         );
  OAI112HS U31283 ( .C1(n27249), .C2(n27257), .A1(n27248), .B1(n27247), .O(
        n13782) );
  OAI112HS U31284 ( .C1(n27258), .C2(n27257), .A1(n27256), .B1(n27255), .O(
        n14168) );
  MUX2S U31285 ( .A(n15889), .B(n27259), .S(gray_img[968]), .O(n27260) );
  AO12S U31286 ( .B1(n15888), .B2(n27261), .A1(n27260), .O(n14125) );
  INV1S U31287 ( .I(gray_img[294]), .O(n27273) );
  INV1S U31288 ( .I(gray_img[292]), .O(n27269) );
  INV1S U31289 ( .I(gray_img[419]), .O(n27266) );
  INV1S U31290 ( .I(gray_img[418]), .O(n27264) );
  INV1S U31291 ( .I(gray_img[417]), .O(n27262) );
  FA1S U31292 ( .A(gray_img[288]), .B(n27262), .CI(gray_img[289]), .CO(n27263)
         );
  FA1S U31293 ( .A(gray_img[290]), .B(n27264), .CI(n27263), .CO(n27265) );
  INV1S U31294 ( .I(n27267), .O(n27268) );
  INV1S U31295 ( .I(gray_img[303]), .O(n27287) );
  INV1S U31296 ( .I(gray_img[302]), .O(n27285) );
  FA1S U31297 ( .A(intadd_16_B_0_), .B(gray_img[425]), .CI(intadd_16_CI), .CO(
        n27276) );
  FA1S U31298 ( .A(n27277), .B(gray_img[426]), .CI(n27276), .CO(n27278) );
  FA1S U31299 ( .A(n27279), .B(gray_img[427]), .CI(n27278), .CO(n27280) );
  FA1S U31300 ( .A(n27281), .B(gray_img[428]), .CI(n27280), .CO(n27282) );
  FA1S U31301 ( .A(n27283), .B(gray_img[429]), .CI(n27282), .CO(n27284) );
  MXL2HS U31302 ( .A(gray_img[302]), .B(gray_img[430]), .S(n30067), .OB(n27301) );
  MXL2HS U31303 ( .A(gray_img[301]), .B(gray_img[429]), .S(n30067), .OB(n27306) );
  MXL2HS U31304 ( .A(gray_img[300]), .B(gray_img[428]), .S(n30067), .OB(n27311) );
  MXL2HS U31305 ( .A(gray_img[299]), .B(gray_img[427]), .S(n30067), .OB(n27317) );
  MXL2HS U31306 ( .A(gray_img[298]), .B(gray_img[426]), .S(n30067), .OB(n27322) );
  MXL2HS U31307 ( .A(gray_img[297]), .B(gray_img[425]), .S(n30067), .OB(n27327) );
  INV1S U31308 ( .I(n27298), .O(n27297) );
  NR2 U31309 ( .I1(n29680), .I2(n27297), .O(n30076) );
  OR2 U31310 ( .I1(n29680), .I2(n27298), .O(n30066) );
  ND2S U31311 ( .I1(n15890), .I2(n30070), .O(n27299) );
  OAI112HS U31312 ( .C1(n30066), .C2(n27301), .A1(n27300), .B1(n27299), .O(
        n27302) );
  ND2S U31313 ( .I1(n26445), .I2(n30070), .O(n27304) );
  OAI112HS U31314 ( .C1(n30066), .C2(n27306), .A1(n27305), .B1(n27304), .O(
        n27307) );
  OAI112HS U31315 ( .C1(n30066), .C2(n27311), .A1(n27310), .B1(n27309), .O(
        n27312) );
  OAI112HS U31316 ( .C1(n30066), .C2(n27317), .A1(n27316), .B1(n27315), .O(
        n27318) );
  OAI112HS U31317 ( .C1(n30066), .C2(n27322), .A1(n27321), .B1(n27320), .O(
        n27323) );
  OAI112HS U31318 ( .C1(n30066), .C2(n27327), .A1(n27326), .B1(n27325), .O(
        n27328) );
  OAI112HS U31319 ( .C1(n27375), .C2(n27332), .A1(n27331), .B1(n27330), .O(
        n27333) );
  MUX2S U31320 ( .A(n30005), .B(n27371), .S(gray_img[20]), .O(n27336) );
  OAI112HS U31321 ( .C1(n27375), .C2(n27337), .A1(n27336), .B1(n27335), .O(
        n27338) );
  OAI112HS U31322 ( .C1(n27375), .C2(n27342), .A1(n27341), .B1(n27340), .O(
        n27343) );
  OAI112HS U31323 ( .C1(n27375), .C2(n27347), .A1(n27346), .B1(n27345), .O(
        n27348) );
  MUX2S U31324 ( .A(gray_img[472]), .B(gray_img[344]), .S(n27353), .O(n27354)
         );
  ND2S U31325 ( .I1(n27355), .I2(n27354), .O(n27360) );
  MUX2S U31326 ( .A(n30005), .B(n27356), .S(gray_img[168]), .O(n27357) );
  OA12S U31327 ( .B1(n29734), .B2(n27358), .A1(n27357), .O(n27359) );
  OAI112HS U31328 ( .C1(n27362), .C2(n27361), .A1(n27360), .B1(n27359), .O(
        n13803) );
  MUX2S U31329 ( .A(gray_img[40]), .B(gray_img[168]), .S(n27363), .O(n27364)
         );
  ND2S U31330 ( .I1(n27365), .I2(n27364), .O(n27368) );
  MUX2S U31331 ( .A(n30005), .B(n27371), .S(gray_img[16]), .O(n27367) );
  ND2S U31332 ( .I1(n15888), .I2(n27371), .O(n27366) );
  ND3S U31333 ( .I1(n27368), .I2(n27367), .I3(n27366), .O(n27369) );
  OAI112HS U31334 ( .C1(n27375), .C2(n27374), .A1(n27373), .B1(n27372), .O(
        n27376) );
  AO12S U31335 ( .B1(n15888), .B2(n27390), .A1(n27383), .O(n14240) );
  INV1S U31336 ( .I(gray_img[236]), .O(n27398) );
  INV1S U31337 ( .I(gray_img[235]), .O(n27396) );
  INV1S U31338 ( .I(gray_img[234]), .O(n27394) );
  INV1S U31339 ( .I(gray_img[233]), .O(n27392) );
  FA1S U31340 ( .A(gray_img[104]), .B(gray_img[105]), .CI(n27392), .CO(n27393)
         );
  FA1S U31341 ( .A(n27394), .B(gray_img[106]), .CI(n27393), .CO(n27395) );
  AOI22S U31342 ( .A1(n27402), .A2(gray_img[237]), .B1(gray_img[238]), .B2(
        n27401), .O(n27403) );
  AOI22S U31343 ( .A1(gray_img[110]), .A2(n27405), .B1(n27404), .B2(n27403), 
        .O(n27408) );
  NR2 U31344 ( .I1(gray_img[111]), .I2(n27406), .O(n27407) );
  INV1S U31345 ( .I(gray_img[103]), .O(n27420) );
  INV1S U31346 ( .I(gray_img[102]), .O(n27418) );
  INV1S U31347 ( .I(gray_img[101]), .O(n27416) );
  INV1S U31348 ( .I(gray_img[99]), .O(n27412) );
  INV1S U31349 ( .I(gray_img[98]), .O(n27410) );
  FA1S U31350 ( .A(gray_img[225]), .B(gray_img[224]), .CI(intadd_125_CI), .CO(
        n27409) );
  FA1S U31351 ( .A(n27410), .B(gray_img[226]), .CI(n27409), .CO(n27411) );
  FA1S U31352 ( .A(n27412), .B(gray_img[227]), .CI(n27411), .CO(n27413) );
  FA1S U31353 ( .A(n27414), .B(gray_img[228]), .CI(n27413), .CO(n27415) );
  FA1S U31354 ( .A(n27416), .B(gray_img[229]), .CI(n27415), .CO(n27417) );
  MXL2HS U31355 ( .A(gray_img[102]), .B(gray_img[230]), .S(n27547), .OB(n27434) );
  MXL2HS U31356 ( .A(gray_img[101]), .B(gray_img[229]), .S(n27547), .OB(n27520) );
  MXL2HS U31357 ( .A(gray_img[100]), .B(gray_img[228]), .S(n27547), .OB(n27525) );
  MXL2HS U31358 ( .A(gray_img[99]), .B(gray_img[227]), .S(n27547), .OB(n27530)
         );
  MXL2HS U31359 ( .A(gray_img[98]), .B(gray_img[226]), .S(n27547), .OB(n27535)
         );
  MXL2HS U31360 ( .A(gray_img[97]), .B(gray_img[225]), .S(n27547), .OB(n27540)
         );
  INV1S U31361 ( .I(n27431), .O(n27430) );
  NR2 U31362 ( .I1(n29680), .I2(n27430), .O(n27556) );
  OR2 U31363 ( .I1(n29680), .I2(n27431), .O(n27546) );
  ND2S U31364 ( .I1(n15890), .I2(n27550), .O(n27432) );
  OAI112HS U31365 ( .C1(n27546), .C2(n27434), .A1(n27433), .B1(n27432), .O(
        n27435) );
  MUX2S U31366 ( .A(n27447), .B(n27446), .S(gray_img[353]), .O(n27441) );
  MUX2S U31367 ( .A(n27447), .B(n27772), .S(gray_img[485]), .O(n27442) );
  MUX2S U31368 ( .A(n27447), .B(n27446), .S(gray_img[352]), .O(n27448) );
  AO12S U31369 ( .B1(n15888), .B2(n27449), .A1(n27448), .O(n14218) );
  INV1S U31370 ( .I(gray_img[365]), .O(n27459) );
  INV1S U31371 ( .I(gray_img[362]), .O(n27453) );
  INV1S U31372 ( .I(gray_img[487]), .O(n27475) );
  INV1S U31373 ( .I(gray_img[486]), .O(n27473) );
  INV1S U31374 ( .I(gray_img[485]), .O(n27471) );
  INV1S U31375 ( .I(gray_img[484]), .O(n27469) );
  INV1S U31376 ( .I(gray_img[483]), .O(n27467) );
  INV1S U31377 ( .I(gray_img[482]), .O(n27465) );
  FA1S U31378 ( .A(gray_img[352]), .B(gray_img[353]), .CI(intadd_115_CI), .CO(
        n27464) );
  FA1S U31379 ( .A(n27465), .B(gray_img[354]), .CI(n27464), .CO(n27466) );
  FA1S U31380 ( .A(n27467), .B(gray_img[355]), .CI(n27466), .CO(n27468) );
  FA1S U31381 ( .A(n27469), .B(gray_img[356]), .CI(n27468), .CO(n27470) );
  FA1S U31382 ( .A(n27471), .B(gray_img[357]), .CI(n27470), .CO(n27472) );
  MXL2HS U31383 ( .A(gray_img[486]), .B(gray_img[358]), .S(n27776), .OB(n27489) );
  MXL2HS U31384 ( .A(gray_img[485]), .B(gray_img[357]), .S(n27776), .OB(n27494) );
  MXL2HS U31385 ( .A(gray_img[484]), .B(gray_img[356]), .S(n27776), .OB(n27499) );
  MXL2HS U31386 ( .A(gray_img[483]), .B(gray_img[355]), .S(n27776), .OB(n27504) );
  MXL2HS U31387 ( .A(gray_img[482]), .B(gray_img[354]), .S(n27776), .OB(n27509) );
  MXL2HS U31388 ( .A(gray_img[481]), .B(gray_img[353]), .S(n27776), .OB(n27515) );
  INV1S U31389 ( .I(n27486), .O(n27485) );
  NR2 U31390 ( .I1(n29680), .I2(n27485), .O(n27785) );
  OR2 U31391 ( .I1(n29680), .I2(n27486), .O(n27775) );
  ND2S U31392 ( .I1(n15890), .I2(n27779), .O(n27487) );
  OAI112HS U31393 ( .C1(n27775), .C2(n27489), .A1(n27488), .B1(n27487), .O(
        n27490) );
  OAI112HS U31394 ( .C1(n27775), .C2(n27494), .A1(n27493), .B1(n27492), .O(
        n27495) );
  OAI112HS U31395 ( .C1(n27775), .C2(n27499), .A1(n27498), .B1(n27497), .O(
        n27500) );
  OAI112HS U31396 ( .C1(n27775), .C2(n27504), .A1(n27503), .B1(n27502), .O(
        n27505) );
  OAI112HS U31397 ( .C1(n27775), .C2(n27509), .A1(n27508), .B1(n27507), .O(
        n27510) );
  OAI112HS U31398 ( .C1(n27775), .C2(n27515), .A1(n27514), .B1(n27513), .O(
        n27516) );
  OAI112HS U31399 ( .C1(n27546), .C2(n27520), .A1(n27519), .B1(n27518), .O(
        n27521) );
  OAI112HS U31400 ( .C1(n27546), .C2(n27525), .A1(n27524), .B1(n27523), .O(
        n27526) );
  OAI112HS U31401 ( .C1(n27546), .C2(n27530), .A1(n27529), .B1(n27528), .O(
        n27531) );
  OAI112HS U31402 ( .C1(n27546), .C2(n27535), .A1(n27534), .B1(n27533), .O(
        n27536) );
  OAI112HS U31403 ( .C1(n27546), .C2(n27540), .A1(n27539), .B1(n27538), .O(
        n27541) );
  AO12S U31404 ( .B1(n15888), .B2(n27545), .A1(n27544), .O(n14262) );
  INV1S U31405 ( .I(n27546), .O(n27549) );
  MUX2S U31406 ( .A(gray_img[96]), .B(gray_img[224]), .S(n27547), .O(n27548)
         );
  ND2S U31407 ( .I1(n27549), .I2(n27548), .O(n27553) );
  MUX2S U31408 ( .A(n29032), .B(n27550), .S(gray_img[48]), .O(n27552) );
  ND2S U31409 ( .I1(n15888), .I2(n27550), .O(n27551) );
  ND3S U31410 ( .I1(n27553), .I2(n27552), .I3(n27551), .O(n27554) );
  FA1S U31411 ( .A(gray_img[121]), .B(gray_img[120]), .CI(intadd_123_CI), .CO(
        n27557) );
  FA1S U31412 ( .A(n27558), .B(gray_img[122]), .CI(n27557), .CO(n27559) );
  FA1S U31413 ( .A(n27560), .B(gray_img[123]), .CI(n27559), .CO(n27561) );
  MXL2HS U31414 ( .A(gray_img[253]), .B(gray_img[125]), .S(n27699), .OB(n27667) );
  INV1S U31415 ( .I(gray_img[246]), .O(n27578) );
  INV1S U31416 ( .I(gray_img[245]), .O(n27576) );
  INV1S U31417 ( .I(gray_img[244]), .O(n27574) );
  INV1S U31418 ( .I(gray_img[243]), .O(n27572) );
  INV1S U31419 ( .I(gray_img[242]), .O(n27570) );
  MXL2HS U31420 ( .A(gray_img[252]), .B(gray_img[124]), .S(n27699), .OB(n27672) );
  MXL2HS U31421 ( .A(gray_img[251]), .B(gray_img[123]), .S(n27699), .OB(n27677) );
  MXL2HS U31422 ( .A(gray_img[250]), .B(gray_img[122]), .S(n27699), .OB(n27682) );
  MUX2S U31423 ( .A(gray_img[241]), .B(gray_img[113]), .S(n27586), .O(n27697)
         );
  MXL2HS U31424 ( .A(gray_img[249]), .B(gray_img[121]), .S(n27699), .OB(n27695) );
  MUX2S U31425 ( .A(gray_img[240]), .B(gray_img[112]), .S(n27586), .O(n27707)
         );
  AOI22S U31426 ( .A1(n27667), .A2(n27669), .B1(n27585), .B2(n27584), .O(
        n27588) );
  MXL2HS U31427 ( .A(gray_img[254]), .B(gray_img[126]), .S(n27699), .OB(n27596) );
  NR2 U31428 ( .I1(n27596), .I2(n27598), .O(n27587) );
  INV1S U31429 ( .I(n27593), .O(n27592) );
  NR2 U31430 ( .I1(n29680), .I2(n27592), .O(n27708) );
  ND2S U31431 ( .I1(n15890), .I2(n27702), .O(n27594) );
  OAI112HS U31432 ( .C1(n27698), .C2(n27596), .A1(n27595), .B1(n27594), .O(
        n27597) );
  INV1S U31433 ( .I(gray_img[503]), .O(n27610) );
  INV1S U31434 ( .I(gray_img[502]), .O(n27608) );
  INV1S U31435 ( .I(gray_img[500]), .O(n27604) );
  INV1S U31436 ( .I(gray_img[499]), .O(n27602) );
  INV1S U31437 ( .I(gray_img[498]), .O(n27600) );
  FA1S U31438 ( .A(gray_img[369]), .B(gray_img[368]), .CI(intadd_112_CI), .CO(
        n27599) );
  FA1S U31439 ( .A(n27600), .B(gray_img[370]), .CI(n27599), .CO(n27601) );
  FA1S U31440 ( .A(n27602), .B(gray_img[371]), .CI(n27601), .CO(n27603) );
  FA1S U31441 ( .A(n27604), .B(gray_img[372]), .CI(n27603), .CO(n27605) );
  FA1S U31442 ( .A(n27606), .B(gray_img[373]), .CI(n27605), .CO(n27607) );
  MXL2HS U31443 ( .A(gray_img[502]), .B(gray_img[374]), .S(n27657), .OB(n27634) );
  INV1S U31444 ( .I(gray_img[509]), .O(n27618) );
  INV1S U31445 ( .I(gray_img[508]), .O(n27616) );
  INV1S U31446 ( .I(gray_img[507]), .O(n27614) );
  INV1S U31447 ( .I(gray_img[506]), .O(n27612) );
  MXL2HS U31448 ( .A(gray_img[501]), .B(gray_img[373]), .S(n27657), .OB(n27639) );
  MXL2HS U31449 ( .A(gray_img[500]), .B(gray_img[372]), .S(n27657), .OB(n27644) );
  MXL2HS U31450 ( .A(gray_img[499]), .B(gray_img[371]), .S(n27657), .OB(n27649) );
  MXL2HS U31451 ( .A(gray_img[498]), .B(gray_img[370]), .S(n27657), .OB(n27654) );
  MUX2S U31452 ( .A(gray_img[505]), .B(gray_img[377]), .S(n27623), .O(n27691)
         );
  MXL2HS U31453 ( .A(gray_img[497]), .B(gray_img[369]), .S(n27657), .OB(n27688) );
  MUX2S U31454 ( .A(gray_img[504]), .B(gray_img[376]), .S(n27623), .O(n27664)
         );
  FA1S U31455 ( .A(n27691), .B(n27688), .CI(n27664), .CO(n27624) );
  INV1S U31456 ( .I(n27631), .O(n27630) );
  NR2 U31457 ( .I1(n29680), .I2(n27630), .O(n27692) );
  OR2 U31458 ( .I1(n29680), .I2(n27631), .O(n27689) );
  ND2S U31459 ( .I1(n15890), .I2(n27685), .O(n27632) );
  OAI112HS U31460 ( .C1(n27689), .C2(n27634), .A1(n27633), .B1(n27632), .O(
        n27635) );
  OAI112HS U31461 ( .C1(n27689), .C2(n27639), .A1(n27638), .B1(n27637), .O(
        n27640) );
  OAI112HS U31462 ( .C1(n27689), .C2(n27644), .A1(n27643), .B1(n27642), .O(
        n27645) );
  OAI112HS U31463 ( .C1(n27689), .C2(n27649), .A1(n27648), .B1(n27647), .O(
        n27650) );
  OAI112HS U31464 ( .C1(n27689), .C2(n27654), .A1(n27653), .B1(n27652), .O(
        n27655) );
  INV1S U31465 ( .I(n27689), .O(n27659) );
  MUX2S U31466 ( .A(gray_img[496]), .B(gray_img[368]), .S(n27657), .O(n27658)
         );
  ND2S U31467 ( .I1(n27659), .I2(n27658), .O(n27662) );
  ND2S U31468 ( .I1(n15888), .I2(n27685), .O(n27660) );
  ND3S U31469 ( .I1(n27662), .I2(n27661), .I3(n27660), .O(n27663) );
  ND2S U31470 ( .I1(n27751), .I2(n27702), .O(n27665) );
  OAI112HS U31471 ( .C1(n27698), .C2(n27667), .A1(n27666), .B1(n27665), .O(
        n27668) );
  OAI112HS U31472 ( .C1(n27698), .C2(n27672), .A1(n27671), .B1(n27670), .O(
        n27673) );
  ND2S U31473 ( .I1(n15887), .I2(n27702), .O(n27675) );
  OAI112HS U31474 ( .C1(n27698), .C2(n27677), .A1(n27676), .B1(n27675), .O(
        n27678) );
  OAI112HS U31475 ( .C1(n27698), .C2(n27682), .A1(n27681), .B1(n27680), .O(
        n27683) );
  OAI112HS U31476 ( .C1(n27689), .C2(n27688), .A1(n27687), .B1(n27686), .O(
        n27690) );
  ND2S U31477 ( .I1(n15928), .I2(n27702), .O(n27693) );
  OAI112HS U31478 ( .C1(n27698), .C2(n27695), .A1(n27694), .B1(n27693), .O(
        n27696) );
  INV1S U31479 ( .I(n27698), .O(n27701) );
  MUX2S U31480 ( .A(gray_img[248]), .B(gray_img[120]), .S(n27699), .O(n27700)
         );
  ND2S U31481 ( .I1(n27701), .I2(n27700), .O(n27705) );
  ND2S U31482 ( .I1(n15888), .I2(n27702), .O(n27703) );
  ND3S U31483 ( .I1(n27705), .I2(n27704), .I3(n27703), .O(n27706) );
  INV1S U31484 ( .I(gray_img[60]), .O(n27715) );
  FA1S U31485 ( .A(gray_img[185]), .B(gray_img[184]), .CI(n27709), .CO(n27710)
         );
  FA1S U31486 ( .A(n27711), .B(gray_img[186]), .CI(n27710), .CO(n27712) );
  FA1S U31487 ( .A(n27713), .B(gray_img[187]), .CI(n27712), .CO(n27714) );
  INV1S U31488 ( .I(gray_img[54]), .O(n27732) );
  INV1S U31489 ( .I(gray_img[53]), .O(n27730) );
  INV1S U31490 ( .I(gray_img[52]), .O(n27728) );
  INV1S U31491 ( .I(gray_img[51]), .O(n27726) );
  INV1S U31492 ( .I(gray_img[50]), .O(n27724) );
  INV1S U31493 ( .I(gray_img[48]), .O(n27722) );
  FA1S U31494 ( .A(intadd_19_B_0_), .B(gray_img[177]), .CI(n27722), .CO(n27723) );
  FA1S U31495 ( .A(n27724), .B(gray_img[178]), .CI(n27723), .CO(n27725) );
  FA1S U31496 ( .A(n27726), .B(gray_img[179]), .CI(n27725), .CO(n27727) );
  FA1S U31497 ( .A(n27728), .B(gray_img[180]), .CI(n27727), .CO(n27729) );
  MAO222 U31498 ( .A1(n27732), .B1(gray_img[182]), .C1(n27731), .O(n27733) );
  MXL2HS U31499 ( .A(gray_img[54]), .B(gray_img[182]), .S(n27786), .OB(n27748)
         );
  MXL2HS U31500 ( .A(gray_img[53]), .B(gray_img[181]), .S(n27786), .OB(n27754)
         );
  MXL2HS U31501 ( .A(gray_img[52]), .B(gray_img[180]), .S(n27786), .OB(n27759)
         );
  MXL2HS U31502 ( .A(gray_img[51]), .B(gray_img[179]), .S(n27786), .OB(n27764)
         );
  MXL2HS U31503 ( .A(gray_img[50]), .B(gray_img[178]), .S(n27786), .OB(n27769)
         );
  MXL2HS U31504 ( .A(gray_img[49]), .B(gray_img[177]), .S(n27786), .OB(n27817)
         );
  MAO222 U31505 ( .A1(n27756), .B1(n27754), .C1(n27739), .O(n27740) );
  MAO222 U31506 ( .A1(n27750), .B1(n27748), .C1(n27740), .O(n27741) );
  INV1S U31507 ( .I(n27745), .O(n27744) );
  NR2 U31508 ( .I1(n29680), .I2(n27744), .O(n27821) );
  OR2 U31509 ( .I1(n29680), .I2(n27745), .O(n27818) );
  ND2S U31510 ( .I1(n15890), .I2(n27814), .O(n27746) );
  OAI112HS U31511 ( .C1(n27818), .C2(n27748), .A1(n27747), .B1(n27746), .O(
        n27749) );
  OAI112HS U31512 ( .C1(n27818), .C2(n27754), .A1(n27753), .B1(n27752), .O(
        n27755) );
  OAI112HS U31513 ( .C1(n27818), .C2(n27759), .A1(n27758), .B1(n27757), .O(
        n27760) );
  OAI112HS U31514 ( .C1(n27818), .C2(n27764), .A1(n27763), .B1(n27762), .O(
        n27765) );
  OAI112HS U31515 ( .C1(n27818), .C2(n27769), .A1(n27768), .B1(n27767), .O(
        n27770) );
  AO12S U31516 ( .B1(n15888), .B2(n27774), .A1(n27773), .O(n14196) );
  INV1S U31517 ( .I(n27775), .O(n27778) );
  MUX2S U31518 ( .A(gray_img[480]), .B(gray_img[352]), .S(n27776), .O(n27777)
         );
  ND2S U31519 ( .I1(n27778), .I2(n27777), .O(n27782) );
  ND2S U31520 ( .I1(n15888), .I2(n27779), .O(n27780) );
  ND3S U31521 ( .I1(n27782), .I2(n27781), .I3(n27780), .O(n27783) );
  INV1S U31522 ( .I(n27818), .O(n27788) );
  MUX2S U31523 ( .A(gray_img[48]), .B(gray_img[176]), .S(n27786), .O(n27787)
         );
  ND2S U31524 ( .I1(n27788), .I2(n27787), .O(n27791) );
  ND2S U31525 ( .I1(n15888), .I2(n27814), .O(n27789) );
  ND3S U31526 ( .I1(n27791), .I2(n27790), .I3(n27789), .O(n27792) );
  MUX2S U31527 ( .A(n15904), .B(n27845), .S(gray_img[157]), .O(n27795) );
  ND2S U31528 ( .I1(n15891), .I2(n27845), .O(n27794) );
  OAI112HS U31529 ( .C1(n27841), .C2(n27796), .A1(n27795), .B1(n27794), .O(
        n27797) );
  OAI112HS U31530 ( .C1(n27841), .C2(n27801), .A1(n27800), .B1(n27799), .O(
        n27802) );
  ND2S U31531 ( .I1(n15887), .I2(n27845), .O(n27804) );
  OAI112HS U31532 ( .C1(n27841), .C2(n27806), .A1(n27805), .B1(n27804), .O(
        n27807) );
  OAI112HS U31533 ( .C1(n27841), .C2(n27811), .A1(n27810), .B1(n27809), .O(
        n27812) );
  OAI112HS U31534 ( .C1(n27818), .C2(n27817), .A1(n27816), .B1(n27815), .O(
        n27819) );
  ND2S U31535 ( .I1(n15928), .I2(n27845), .O(n27822) );
  OAI112HS U31536 ( .C1(n27841), .C2(n27824), .A1(n27823), .B1(n27822), .O(
        n27825) );
  AO12S U31537 ( .B1(n15888), .B2(n27829), .A1(n27828), .O(n14108) );
  INV1S U31538 ( .I(n27830), .O(n27833) );
  MUX2S U31539 ( .A(gray_img[992]), .B(gray_img[864]), .S(n27831), .O(n27832)
         );
  ND2S U31540 ( .I1(n27833), .I2(n27832), .O(n27837) );
  ND2S U31541 ( .I1(n15888), .I2(n27834), .O(n27835) );
  ND3S U31542 ( .I1(n27837), .I2(n27836), .I3(n27835), .O(n27838) );
  INV1S U31543 ( .I(n27841), .O(n27844) );
  MUX2S U31544 ( .A(gray_img[304]), .B(gray_img[432]), .S(n27842), .O(n27843)
         );
  ND2S U31545 ( .I1(n27844), .I2(n27843), .O(n27848) );
  ND2S U31546 ( .I1(n15888), .I2(n27845), .O(n27846) );
  ND3S U31547 ( .I1(n27848), .I2(n27847), .I3(n27846), .O(n27849) );
  INV1S U31548 ( .I(gray_img[21]), .O(n27859) );
  INV1S U31549 ( .I(gray_img[20]), .O(n27857) );
  INV1S U31550 ( .I(gray_img[18]), .O(n27853) );
  FA1S U31551 ( .A(intadd_11_B_0_), .B(gray_img[145]), .CI(intadd_11_CI), .CO(
        n27852) );
  FA1S U31552 ( .A(n27853), .B(gray_img[146]), .CI(n27852), .CO(n27854) );
  FA1S U31553 ( .A(n27855), .B(gray_img[147]), .CI(n27854), .CO(n27856) );
  FA1S U31554 ( .A(n27857), .B(gray_img[148]), .CI(n27856), .CO(n27858) );
  MXL2HS U31555 ( .A(gray_img[22]), .B(gray_img[150]), .S(n30078), .OB(n27892)
         );
  INV1S U31556 ( .I(gray_img[154]), .O(n27866) );
  FA1S U31557 ( .A(gray_img[25]), .B(gray_img[24]), .CI(n27864), .CO(n27865)
         );
  FA1S U31558 ( .A(n27866), .B(gray_img[26]), .CI(n27865), .CO(n27867) );
  FA1S U31559 ( .A(n27868), .B(gray_img[27]), .CI(n27867), .CO(n27869) );
  MXL2HS U31560 ( .A(gray_img[21]), .B(gray_img[149]), .S(n30078), .OB(n28822)
         );
  MXL2HS U31561 ( .A(gray_img[20]), .B(gray_img[148]), .S(n30078), .OB(n28827)
         );
  MXL2HS U31562 ( .A(gray_img[19]), .B(gray_img[147]), .S(n30078), .OB(n28832)
         );
  MXL2HS U31563 ( .A(gray_img[18]), .B(gray_img[146]), .S(n30078), .OB(n28837)
         );
  MXL2HS U31564 ( .A(gray_img[17]), .B(gray_img[145]), .S(n30078), .OB(n28850)
         );
  OR2 U31565 ( .I1(n29680), .I2(n27886), .O(n30077) );
  INV1S U31566 ( .I(n27886), .O(n27887) );
  OA12S U31567 ( .B1(gray_img[14]), .B2(n29427), .A1(n30081), .O(n27889) );
  MOAI1S U31568 ( .A1(n30081), .A2(gray_img[14]), .B1(n29825), .B2(n27889), 
        .O(n27890) );
  OAI112HS U31569 ( .C1(n27892), .C2(n30077), .A1(n27891), .B1(n27890), .O(
        n13748) );
  INV1S U31570 ( .I(gray_img[1535]), .O(n27904) );
  INV1S U31571 ( .I(gray_img[1534]), .O(n27902) );
  INV1S U31572 ( .I(gray_img[1533]), .O(n27900) );
  INV1S U31573 ( .I(gray_img[1530]), .O(n27894) );
  MXL2HS U31574 ( .A(gray_img[1534]), .B(gray_img[1406]), .S(n27918), .OB(
        n27933) );
  INV1S U31575 ( .I(gray_img[1396]), .O(n27911) );
  FA1S U31576 ( .A(gray_img[1521]), .B(gray_img[1520]), .CI(n27905), .CO(
        n27906) );
  FA1S U31577 ( .A(n27907), .B(gray_img[1522]), .CI(n27906), .CO(n27908) );
  FA1S U31578 ( .A(n27909), .B(gray_img[1523]), .CI(n27908), .CO(n27910) );
  MXL2HS U31579 ( .A(gray_img[1533]), .B(gray_img[1405]), .S(n27918), .OB(
        n27938) );
  MXL2HS U31580 ( .A(gray_img[1532]), .B(gray_img[1404]), .S(n27918), .OB(
        n27943) );
  MXL2HS U31581 ( .A(gray_img[1531]), .B(gray_img[1403]), .S(n27918), .OB(
        n27948) );
  MXL2HS U31582 ( .A(gray_img[1530]), .B(gray_img[1402]), .S(n27918), .OB(
        n27953) );
  MXL2HS U31583 ( .A(gray_img[1528]), .B(gray_img[1400]), .S(n27918), .OB(
        n28143) );
  MXL2HS U31584 ( .A(gray_img[1529]), .B(gray_img[1401]), .S(n27918), .OB(
        n27958) );
  INV1S U31585 ( .I(n28137), .O(n28139) );
  OAI112HS U31586 ( .C1(n27933), .C2(n28142), .A1(n27932), .B1(n27931), .O(
        n13925) );
  OAI112HS U31587 ( .C1(n27938), .C2(n28142), .A1(n27937), .B1(n27936), .O(
        n13926) );
  OAI112HS U31588 ( .C1(n27943), .C2(n28142), .A1(n27942), .B1(n27941), .O(
        n13927) );
  OAI112HS U31589 ( .C1(n27948), .C2(n28142), .A1(n27947), .B1(n27946), .O(
        n14671) );
  OAI112HS U31590 ( .C1(n27953), .C2(n28142), .A1(n27952), .B1(n27951), .O(
        n13672) );
  OAI112HS U31591 ( .C1(n27958), .C2(n28142), .A1(n27957), .B1(n27956), .O(
        n13696) );
  ND2S U31592 ( .I1(n28201), .I2(gray_img[1381]), .O(n27960) );
  INV1S U31593 ( .I(gray_img[1381]), .O(n27993) );
  OAI112HS U31594 ( .C1(n29831), .C2(n28201), .A1(n27960), .B1(n27959), .O(
        n15160) );
  INV1S U31595 ( .I(n28201), .O(n28203) );
  MUX2S U31596 ( .A(n15889), .B(n27969), .S(gray_img[1506]), .O(n27964) );
  MUX2S U31597 ( .A(n27447), .B(n27969), .S(gray_img[1504]), .O(n27965) );
  AO12S U31598 ( .B1(n15888), .B2(n27971), .A1(n27965), .O(n13936) );
  MUX2S U31599 ( .A(n15889), .B(n27969), .S(gray_img[1505]), .O(n27970) );
  INV1S U31600 ( .I(gray_img[1518]), .O(n27982) );
  INV1S U31601 ( .I(gray_img[1517]), .O(n27980) );
  INV1S U31602 ( .I(gray_img[1516]), .O(n27978) );
  INV1S U31603 ( .I(gray_img[1515]), .O(n27976) );
  INV1S U31604 ( .I(gray_img[1514]), .O(n27974) );
  FA1S U31605 ( .A(gray_img[1385]), .B(gray_img[1384]), .CI(intadd_55_CI), 
        .CO(n27973) );
  FA1S U31606 ( .A(n27974), .B(gray_img[1386]), .CI(n27973), .CO(n27975) );
  FA1S U31607 ( .A(n27976), .B(gray_img[1387]), .CI(n27975), .CO(n27977) );
  FA1S U31608 ( .A(n27978), .B(gray_img[1388]), .CI(n27977), .CO(n27979) );
  INV1S U31609 ( .I(gray_img[1506]), .O(n27988) );
  INV1S U31610 ( .I(gray_img[1505]), .O(n27986) );
  FA1S U31611 ( .A(n27986), .B(n27985), .CI(gray_img[1377]), .CO(n27987) );
  FA1S U31612 ( .A(gray_img[1378]), .B(n27988), .CI(n27987), .CO(n27989) );
  FA1S U31613 ( .A(gray_img[1379]), .B(n27990), .CI(n27989), .CO(n27991) );
  NR2 U31614 ( .I1(gray_img[1509]), .I2(n27993), .O(n27994) );
  MOAI1S U31615 ( .A1(n27995), .A2(n27994), .B1(gray_img[1509]), .B2(n27993), 
        .O(n27996) );
  OAI12HS U31616 ( .B1(gray_img[1510]), .B2(n27997), .A1(n27996), .O(n28000)
         );
  ND2S U31617 ( .I1(n28002), .I2(gray_img[1511]), .O(n27999) );
  ND2S U31618 ( .I1(n27997), .I2(gray_img[1510]), .O(n27998) );
  OAI12HS U31619 ( .B1(gray_img[1511]), .B2(n28002), .A1(n28001), .O(n28205)
         );
  MXL2HS U31620 ( .A(gray_img[1510]), .B(gray_img[1382]), .S(n28205), .OB(
        n28016) );
  MXL2HS U31621 ( .A(gray_img[1509]), .B(gray_img[1381]), .S(n28205), .OB(
        n28103) );
  MXL2HS U31622 ( .A(gray_img[1508]), .B(gray_img[1380]), .S(n28205), .OB(
        n28108) );
  MXL2HS U31623 ( .A(gray_img[1507]), .B(gray_img[1379]), .S(n28205), .OB(
        n28113) );
  MXL2HS U31624 ( .A(gray_img[1506]), .B(gray_img[1378]), .S(n28205), .OB(
        n28118) );
  MXL2HS U31625 ( .A(gray_img[1505]), .B(gray_img[1377]), .S(n28205), .OB(
        n28131) );
  INV1S U31626 ( .I(n28013), .O(n28012) );
  NR2 U31627 ( .I1(n29680), .I2(n28012), .O(n28214) );
  OR2 U31628 ( .I1(n29680), .I2(n28013), .O(n28204) );
  ND2S U31629 ( .I1(n15890), .I2(n28208), .O(n28014) );
  OAI112HS U31630 ( .C1(n28204), .C2(n28016), .A1(n28015), .B1(n28014), .O(
        n28017) );
  MUX2S U31631 ( .A(n27447), .B(n28090), .S(gray_img[1121]), .O(n28023) );
  MUX2S U31632 ( .A(n15889), .B(n28029), .S(gray_img[1252]), .O(n28025) );
  MUX2S U31633 ( .A(n15889), .B(n28029), .S(gray_img[1251]), .O(n28026) );
  MUX2S U31634 ( .A(n15889), .B(n28029), .S(gray_img[1250]), .O(n28027) );
  MUX2S U31635 ( .A(n27447), .B(n28029), .S(gray_img[1248]), .O(n28028) );
  AO12S U31636 ( .B1(n19092), .B2(n28031), .A1(n28028), .O(n14020) );
  MUX2S U31637 ( .A(n15889), .B(n28029), .S(gray_img[1249]), .O(n28030) );
  INV1S U31638 ( .I(gray_img[1252]), .O(n28037) );
  INV1S U31639 ( .I(gray_img[1251]), .O(n28035) );
  INV1S U31640 ( .I(gray_img[1250]), .O(n28033) );
  FA1S U31641 ( .A(intadd_72_B_0_), .B(gray_img[1121]), .CI(intadd_72_CI), 
        .CO(n28032) );
  FA1S U31642 ( .A(n28033), .B(gray_img[1122]), .CI(n28032), .CO(n28034) );
  FA1S U31643 ( .A(n28035), .B(gray_img[1123]), .CI(n28034), .CO(n28036) );
  MXL2HS U31644 ( .A(gray_img[1254]), .B(gray_img[1126]), .S(n28093), .OB(
        n28067) );
  INV1S U31645 ( .I(gray_img[1132]), .O(n28049) );
  MXL2HS U31646 ( .A(gray_img[1253]), .B(gray_img[1125]), .S(n28093), .OB(
        n28072) );
  MXL2HS U31647 ( .A(gray_img[1252]), .B(gray_img[1124]), .S(n28093), .OB(
        n28077) );
  MXL2HS U31648 ( .A(gray_img[1251]), .B(gray_img[1123]), .S(n28093), .OB(
        n28082) );
  MUX2S U31649 ( .A(gray_img[1130]), .B(gray_img[1258]), .S(n28056), .O(n28089) );
  MXL2HS U31650 ( .A(gray_img[1250]), .B(gray_img[1122]), .S(n28093), .OB(
        n28087) );
  MUX2S U31651 ( .A(gray_img[1128]), .B(gray_img[1256]), .S(n28056), .O(n28100) );
  MXL2HS U31652 ( .A(gray_img[1249]), .B(gray_img[1121]), .S(n28093), .OB(
        n28124) );
  MUX2S U31653 ( .A(gray_img[1129]), .B(gray_img[1257]), .S(n28056), .O(n28127) );
  FA1S U31654 ( .A(n28100), .B(n28124), .CI(n28127), .CO(n28057) );
  INV1S U31655 ( .I(n28064), .O(n28063) );
  NR2 U31656 ( .I1(n29680), .I2(n28063), .O(n28128) );
  OR2 U31657 ( .I1(n29680), .I2(n28064), .O(n28125) );
  ND2S U31658 ( .I1(n15890), .I2(n28121), .O(n28065) );
  OAI112HS U31659 ( .C1(n28125), .C2(n28067), .A1(n28066), .B1(n28065), .O(
        n28068) );
  ND2S U31660 ( .I1(n26828), .I2(n28121), .O(n28070) );
  OAI112HS U31661 ( .C1(n28125), .C2(n28072), .A1(n28071), .B1(n28070), .O(
        n28073) );
  OAI112HS U31662 ( .C1(n28125), .C2(n28077), .A1(n28076), .B1(n28075), .O(
        n28078) );
  OAI112HS U31663 ( .C1(n28125), .C2(n28082), .A1(n28081), .B1(n28080), .O(
        n28083) );
  OAI112HS U31664 ( .C1(n28125), .C2(n28087), .A1(n28086), .B1(n28085), .O(
        n28088) );
  AO12S U31665 ( .B1(n15888), .B2(n28092), .A1(n28091), .O(n14078) );
  INV1S U31666 ( .I(n28125), .O(n28095) );
  MUX2S U31667 ( .A(gray_img[1248]), .B(gray_img[1120]), .S(n28093), .O(n28094) );
  ND2S U31668 ( .I1(n28095), .I2(n28094), .O(n28098) );
  ND2S U31669 ( .I1(n15888), .I2(n28121), .O(n28096) );
  ND3S U31670 ( .I1(n28098), .I2(n28097), .I3(n28096), .O(n28099) );
  ND2S U31671 ( .I1(n26445), .I2(n28208), .O(n28101) );
  OAI112HS U31672 ( .C1(n28204), .C2(n28103), .A1(n28102), .B1(n28101), .O(
        n28104) );
  OAI112HS U31673 ( .C1(n28204), .C2(n28108), .A1(n28107), .B1(n28106), .O(
        n28109) );
  OAI112HS U31674 ( .C1(n28204), .C2(n28113), .A1(n28112), .B1(n28111), .O(
        n28114) );
  OAI112HS U31675 ( .C1(n28204), .C2(n28118), .A1(n28117), .B1(n28116), .O(
        n28119) );
  OAI112HS U31676 ( .C1(n28125), .C2(n28124), .A1(n28123), .B1(n28122), .O(
        n28126) );
  OAI112HS U31677 ( .C1(n28204), .C2(n28131), .A1(n28130), .B1(n28129), .O(
        n28132) );
  MUX2S U31678 ( .A(gray_img[1392]), .B(gray_img[1520]), .S(n28134), .O(n28135) );
  OAI112HS U31679 ( .C1(n28143), .C2(n28142), .A1(n28141), .B1(n28140), .O(
        n13723) );
  INV1S U31680 ( .I(gray_img[573]), .O(n28151) );
  MAO222S U31681 ( .A1(intadd_189_B_0_), .B1(intadd_189_A_0_), .C1(
        gray_img[697]), .O(n28144) );
  FA1S U31682 ( .A(gray_img[698]), .B(n28145), .CI(n28144), .CO(n28146) );
  FA1S U31683 ( .A(gray_img[699]), .B(n28147), .CI(n28146), .CO(n28148) );
  FA1S U31684 ( .A(gray_img[700]), .B(n28149), .CI(n28148), .CO(n28150) );
  FA1S U31685 ( .A(gray_img[701]), .B(n28151), .CI(n28150), .CO(n28152) );
  NR2 U31686 ( .I1(n28154), .I2(n28155), .O(n28157) );
  AOI12HS U31687 ( .B1(n28155), .B2(n28154), .A1(gray_img[703]), .O(n28156) );
  MXL2HS U31688 ( .A(gray_img[574]), .B(gray_img[702]), .S(n28170), .OB(n28185) );
  INV1S U31689 ( .I(gray_img[694]), .O(n28167) );
  INV1S U31690 ( .I(gray_img[693]), .O(n28165) );
  INV1S U31691 ( .I(gray_img[692]), .O(n28163) );
  INV1S U31692 ( .I(gray_img[691]), .O(n28161) );
  INV1S U31693 ( .I(gray_img[690]), .O(n28159) );
  FA1S U31694 ( .A(gray_img[561]), .B(gray_img[560]), .CI(intadd_142_CI), .CO(
        n28158) );
  FA1S U31695 ( .A(n28159), .B(gray_img[562]), .CI(n28158), .CO(n28160) );
  FA1S U31696 ( .A(n28161), .B(gray_img[563]), .CI(n28160), .CO(n28162) );
  FA1S U31697 ( .A(n28163), .B(gray_img[564]), .CI(n28162), .CO(n28164) );
  MXL2HS U31698 ( .A(gray_img[573]), .B(gray_img[701]), .S(n28170), .OB(n28254) );
  MXL2HS U31699 ( .A(gray_img[572]), .B(gray_img[700]), .S(n28170), .OB(n28190) );
  MXL2HS U31700 ( .A(gray_img[571]), .B(gray_img[699]), .S(n28170), .OB(n28195) );
  MXL2HS U31701 ( .A(gray_img[570]), .B(gray_img[698]), .S(n28170), .OB(n28200) );
  MXL2HS U31702 ( .A(gray_img[568]), .B(gray_img[696]), .S(n28170), .OB(n28220) );
  MXL2HS U31703 ( .A(gray_img[569]), .B(gray_img[697]), .S(n28170), .OB(n28240) );
  OR2 U31704 ( .I1(n29680), .I2(n28179), .O(n28253) );
  INV1S U31705 ( .I(n28179), .O(n28180) );
  INV1S U31706 ( .I(n28248), .O(n28250) );
  OAI112HS U31707 ( .C1(n28185), .C2(n28253), .A1(n28184), .B1(n28183), .O(
        n13652) );
  OAI112HS U31708 ( .C1(n28190), .C2(n28253), .A1(n28189), .B1(n28188), .O(
        n13654) );
  OAI112HS U31709 ( .C1(n28195), .C2(n28253), .A1(n28194), .B1(n28193), .O(
        n13655) );
  OAI112HS U31710 ( .C1(n28200), .C2(n28253), .A1(n28199), .B1(n28198), .O(
        n14670) );
  INV1S U31711 ( .I(n28204), .O(n28207) );
  MUX2S U31712 ( .A(gray_img[1504]), .B(gray_img[1376]), .S(n28205), .O(n28206) );
  ND2S U31713 ( .I1(n28207), .I2(n28206), .O(n28211) );
  ND2S U31714 ( .I1(n15888), .I2(n28208), .O(n28209) );
  ND3S U31715 ( .I1(n28211), .I2(n28210), .I3(n28209), .O(n28212) );
  MUX2S U31716 ( .A(gray_img[688]), .B(gray_img[560]), .S(n28215), .O(n28216)
         );
  OAI112HS U31717 ( .C1(n28220), .C2(n28253), .A1(n28219), .B1(n28218), .O(
        n13783) );
  INV1S U31718 ( .I(n28728), .O(n28730) );
  OAI112HS U31719 ( .C1(n28225), .C2(n28733), .A1(n28224), .B1(n28223), .O(
        n14872) );
  OAI112HS U31720 ( .C1(n28230), .C2(n28733), .A1(n28229), .B1(n28228), .O(
        n14672) );
  OAI112HS U31721 ( .C1(n28235), .C2(n28733), .A1(n28234), .B1(n28233), .O(
        n14471) );
  OAI112HS U31722 ( .C1(n28240), .C2(n28253), .A1(n28239), .B1(n28238), .O(
        n14273) );
  OAI112HS U31723 ( .C1(n28245), .C2(n28733), .A1(n28244), .B1(n28243), .O(
        n14269) );
  OAI112HS U31724 ( .C1(n28254), .C2(n28253), .A1(n28252), .B1(n28251), .O(
        n13653) );
  OAI112HS U31725 ( .C1(n28259), .C2(n28733), .A1(n28258), .B1(n28257), .O(
        n15074) );
  MUX2S U31726 ( .A(n15889), .B(n28269), .S(gray_img[1237]), .O(n28260) );
  MUX2S U31727 ( .A(n15889), .B(n28269), .S(gray_img[1235]), .O(n28262) );
  MUX2S U31728 ( .A(n15889), .B(n28269), .S(gray_img[1234]), .O(n28263) );
  MUX2S U31729 ( .A(n15889), .B(n28269), .S(gray_img[1232]), .O(n28264) );
  AO12S U31730 ( .B1(n19092), .B2(n28271), .A1(n28264), .O(n14029) );
  MUX2S U31731 ( .A(n15889), .B(n28421), .S(gray_img[1108]), .O(n28266) );
  MUX2S U31732 ( .A(n15889), .B(n28421), .S(gray_img[1107]), .O(n28267) );
  MUX2S U31733 ( .A(n15889), .B(n28421), .S(gray_img[1106]), .O(n28268) );
  MUX2S U31734 ( .A(n15889), .B(n28269), .S(gray_img[1233]), .O(n28270) );
  MUX2S U31735 ( .A(n15889), .B(n28421), .S(gray_img[1105]), .O(n28272) );
  MUX2S U31736 ( .A(n27447), .B(n28282), .S(gray_img[1117]), .O(n28273) );
  MUX2S U31737 ( .A(n15889), .B(n28282), .S(gray_img[1115]), .O(n28275) );
  MUX2S U31738 ( .A(n15889), .B(n28282), .S(gray_img[1114]), .O(n28276) );
  MUX2S U31739 ( .A(n15889), .B(n28282), .S(gray_img[1113]), .O(n28277) );
  MUX2S U31740 ( .A(n15889), .B(n28286), .S(gray_img[1244]), .O(n28279) );
  MUX2S U31741 ( .A(n15889), .B(n28286), .S(gray_img[1243]), .O(n28280) );
  MUX2S U31742 ( .A(n15889), .B(n28286), .S(gray_img[1242]), .O(n28281) );
  AO12S U31743 ( .B1(n19092), .B2(n28284), .A1(n28283), .O(n14079) );
  MUX2S U31744 ( .A(n15889), .B(n28286), .S(gray_img[1241]), .O(n28285) );
  MUX2S U31745 ( .A(n15889), .B(n28286), .S(gray_img[1240]), .O(n28287) );
  AO12S U31746 ( .B1(n19092), .B2(n28288), .A1(n28287), .O(n14028) );
  INV1S U31747 ( .I(gray_img[1246]), .O(n28299) );
  INV1S U31748 ( .I(gray_img[1245]), .O(n28297) );
  INV1S U31749 ( .I(gray_img[1244]), .O(n28295) );
  INV1S U31750 ( .I(gray_img[1243]), .O(n28293) );
  INV1S U31751 ( .I(gray_img[1242]), .O(n28291) );
  FA1S U31752 ( .A(gray_img[1112]), .B(gray_img[1113]), .CI(n28289), .CO(
        n28290) );
  FA1S U31753 ( .A(n28291), .B(gray_img[1114]), .CI(n28290), .CO(n28292) );
  FA1S U31754 ( .A(n28293), .B(gray_img[1115]), .CI(n28292), .CO(n28294) );
  FA1S U31755 ( .A(n28295), .B(gray_img[1116]), .CI(n28294), .CO(n28296) );
  INV1S U31756 ( .I(gray_img[1111]), .O(n28314) );
  INV1S U31757 ( .I(gray_img[1110]), .O(n28312) );
  INV1S U31758 ( .I(gray_img[1109]), .O(n28310) );
  INV1S U31759 ( .I(gray_img[1108]), .O(n28308) );
  INV1S U31760 ( .I(gray_img[1107]), .O(n28306) );
  INV1S U31761 ( .I(gray_img[1106]), .O(n28304) );
  INV1S U31762 ( .I(gray_img[1105]), .O(n28302) );
  FA1S U31763 ( .A(n28308), .B(gray_img[1236]), .CI(n28307), .CO(n28309) );
  FA1S U31764 ( .A(n28310), .B(gray_img[1237]), .CI(n28309), .CO(n28311) );
  MXL2HS U31765 ( .A(gray_img[1110]), .B(gray_img[1238]), .S(n28424), .OB(
        n28328) );
  MXL2HS U31766 ( .A(gray_img[1109]), .B(gray_img[1237]), .S(n28424), .OB(
        n28403) );
  MXL2HS U31767 ( .A(gray_img[1108]), .B(gray_img[1236]), .S(n28424), .OB(
        n28408) );
  MXL2HS U31768 ( .A(gray_img[1107]), .B(gray_img[1235]), .S(n28424), .OB(
        n28413) );
  MXL2HS U31769 ( .A(gray_img[1106]), .B(gray_img[1234]), .S(n28424), .OB(
        n28418) );
  MXL2HS U31770 ( .A(gray_img[1105]), .B(gray_img[1233]), .S(n28424), .OB(
        n28455) );
  INV1S U31771 ( .I(n28325), .O(n28324) );
  NR2 U31772 ( .I1(n29680), .I2(n28324), .O(n28459) );
  ND2S U31773 ( .I1(n15890), .I2(n28452), .O(n28326) );
  OAI112HS U31774 ( .C1(n28456), .C2(n28328), .A1(n28327), .B1(n28326), .O(
        n28329) );
  MUX2S U31775 ( .A(n27447), .B(n28594), .S(gray_img[1363]), .O(n28338) );
  MUX2S U31776 ( .A(n15889), .B(n28594), .S(gray_img[1362]), .O(n28339) );
  MUX2S U31777 ( .A(n15889), .B(n28353), .S(gray_img[1500]), .O(n28345) );
  MUX2S U31778 ( .A(n15889), .B(n28353), .S(gray_img[1499]), .O(n28346) );
  MUX2S U31779 ( .A(n27447), .B(n28353), .S(gray_img[1496]), .O(n28348) );
  AO12S U31780 ( .B1(n19092), .B2(n28355), .A1(n28348), .O(n13942) );
  MUX2S U31781 ( .A(n15889), .B(n28357), .S(gray_img[1371]), .O(n28351) );
  MUX2S U31782 ( .A(n15889), .B(n28357), .S(gray_img[1370]), .O(n28352) );
  MUX2S U31783 ( .A(n15889), .B(n28353), .S(gray_img[1497]), .O(n28354) );
  MUX2S U31784 ( .A(n27447), .B(n28357), .S(gray_img[1369]), .O(n28356) );
  MUX2S U31785 ( .A(n15889), .B(n28357), .S(gray_img[1368]), .O(n28358) );
  AO12S U31786 ( .B1(n19092), .B2(n28359), .A1(n28358), .O(n13991) );
  INV1S U31787 ( .I(gray_img[1373]), .O(n28368) );
  INV1S U31788 ( .I(gray_img[1372]), .O(n28366) );
  INV1S U31789 ( .I(gray_img[1370]), .O(n28362) );
  FA1S U31790 ( .A(n28362), .B(gray_img[1498]), .CI(n28361), .CO(n28363) );
  FA1S U31791 ( .A(n28364), .B(gray_img[1499]), .CI(n28363), .CO(n28365) );
  FA1S U31792 ( .A(n28366), .B(gray_img[1500]), .CI(n28365), .CO(n28367) );
  INV1S U31793 ( .I(gray_img[1367]), .O(n28384) );
  INV1S U31794 ( .I(gray_img[1366]), .O(n28382) );
  FA1S U31795 ( .A(gray_img[1489]), .B(gray_img[1488]), .CI(intadd_140_CI), 
        .CO(n28373) );
  FA1S U31796 ( .A(n28374), .B(gray_img[1490]), .CI(n28373), .CO(n28375) );
  FA1S U31797 ( .A(n28376), .B(gray_img[1491]), .CI(n28375), .CO(n28377) );
  FA1S U31798 ( .A(n28378), .B(gray_img[1492]), .CI(n28377), .CO(n28379) );
  FA1S U31799 ( .A(n28380), .B(gray_img[1493]), .CI(n28379), .CO(n28381) );
  MXL2HS U31800 ( .A(gray_img[1366]), .B(gray_img[1494]), .S(n28598), .OB(
        n28398) );
  MXL2HS U31801 ( .A(gray_img[1365]), .B(gray_img[1493]), .S(n28598), .OB(
        n28434) );
  MXL2HS U31802 ( .A(gray_img[1364]), .B(gray_img[1492]), .S(n28598), .OB(
        n28439) );
  MXL2HS U31803 ( .A(gray_img[1363]), .B(gray_img[1491]), .S(n28598), .OB(
        n28444) );
  MXL2HS U31804 ( .A(gray_img[1362]), .B(gray_img[1490]), .S(n28598), .OB(
        n28449) );
  MUX2S U31805 ( .A(gray_img[1369]), .B(gray_img[1497]), .S(n28385), .O(n28464) );
  MXL2HS U31806 ( .A(gray_img[1361]), .B(gray_img[1489]), .S(n28598), .OB(
        n28462) );
  INV1S U31807 ( .I(n28395), .O(n28394) );
  NR2 U31808 ( .I1(n29680), .I2(n28394), .O(n28607) );
  MUX2S U31809 ( .A(n15904), .B(n28601), .S(gray_img[686]), .O(n28397) );
  ND2S U31810 ( .I1(n15890), .I2(n28601), .O(n28396) );
  OAI112HS U31811 ( .C1(n28597), .C2(n28398), .A1(n28397), .B1(n28396), .O(
        n28399) );
  ND2S U31812 ( .I1(n27751), .I2(n28452), .O(n28401) );
  OAI112HS U31813 ( .C1(n28456), .C2(n28403), .A1(n28402), .B1(n28401), .O(
        n28404) );
  OAI112HS U31814 ( .C1(n28456), .C2(n28408), .A1(n28407), .B1(n28406), .O(
        n28409) );
  OAI112HS U31815 ( .C1(n28456), .C2(n28413), .A1(n28412), .B1(n28411), .O(
        n28414) );
  OAI112HS U31816 ( .C1(n28456), .C2(n28418), .A1(n28417), .B1(n28416), .O(
        n28419) );
  MUX2S U31817 ( .A(n15889), .B(n28421), .S(gray_img[1104]), .O(n28422) );
  AO12S U31818 ( .B1(n15888), .B2(n28423), .A1(n28422), .O(n14080) );
  INV1S U31819 ( .I(n28456), .O(n28426) );
  MUX2S U31820 ( .A(gray_img[1104]), .B(gray_img[1232]), .S(n28424), .O(n28425) );
  ND2S U31821 ( .I1(n28426), .I2(n28425), .O(n28429) );
  MUX2S U31822 ( .A(n29032), .B(n28452), .S(gray_img[552]), .O(n28428) );
  ND2S U31823 ( .I1(n15888), .I2(n28452), .O(n28427) );
  ND3S U31824 ( .I1(n28429), .I2(n28428), .I3(n28427), .O(n28430) );
  MUX2S U31825 ( .A(n15904), .B(n28601), .S(gray_img[685]), .O(n28433) );
  ND2S U31826 ( .I1(n26828), .I2(n28601), .O(n28432) );
  OAI112HS U31827 ( .C1(n28597), .C2(n28434), .A1(n28433), .B1(n28432), .O(
        n28435) );
  OAI112HS U31828 ( .C1(n28597), .C2(n28439), .A1(n28438), .B1(n28437), .O(
        n28440) );
  OAI112HS U31829 ( .C1(n28597), .C2(n28444), .A1(n28443), .B1(n28442), .O(
        n28445) );
  OAI112HS U31830 ( .C1(n28597), .C2(n28449), .A1(n28448), .B1(n28447), .O(
        n28450) );
  OAI112HS U31831 ( .C1(n28456), .C2(n28455), .A1(n28454), .B1(n28453), .O(
        n28457) );
  OAI112HS U31832 ( .C1(n28597), .C2(n28462), .A1(n28461), .B1(n28460), .O(
        n28463) );
  MUX2S U31833 ( .A(n15889), .B(n28473), .S(gray_img[1228]), .O(n28466) );
  MUX2S U31834 ( .A(n15889), .B(n28473), .S(gray_img[1227]), .O(n28468) );
  MUX2S U31835 ( .A(n15889), .B(n28473), .S(gray_img[1226]), .O(n28469) );
  MUX2S U31836 ( .A(n27447), .B(n28473), .S(gray_img[1224]), .O(n28470) );
  AO12S U31837 ( .B1(n15888), .B2(n28475), .A1(n28470), .O(n14037) );
  MUX2S U31838 ( .A(n15889), .B(n28478), .S(gray_img[1099]), .O(n28471) );
  MUX2S U31839 ( .A(n15889), .B(n28478), .S(gray_img[1098]), .O(n28472) );
  MUX2S U31840 ( .A(n27447), .B(n28473), .S(gray_img[1225]), .O(n28474) );
  MUX2S U31841 ( .A(n15889), .B(n28478), .S(gray_img[1097]), .O(n28476) );
  MUX2S U31842 ( .A(n15889), .B(n28478), .S(gray_img[1100]), .O(n28477) );
  MUX2S U31843 ( .A(n15889), .B(n28478), .S(gray_img[1096]), .O(n28479) );
  AO12S U31844 ( .B1(n15888), .B2(n28480), .A1(n28479), .O(n14081) );
  INV1S U31845 ( .I(gray_img[1231]), .O(n28494) );
  INV1S U31846 ( .I(gray_img[1230]), .O(n28492) );
  INV1S U31847 ( .I(gray_img[1229]), .O(n28490) );
  INV1S U31848 ( .I(gray_img[1099]), .O(n28485) );
  INV1S U31849 ( .I(gray_img[1097]), .O(n28481) );
  FA1S U31850 ( .A(gray_img[1225]), .B(gray_img[1224]), .CI(n28481), .CO(
        n28482) );
  INV1S U31851 ( .I(n28486), .O(n28488) );
  INV1S U31852 ( .I(gray_img[1228]), .O(n28487) );
  FA1S U31853 ( .A(n28488), .B(n28487), .CI(gray_img[1100]), .CO(n28489) );
  FA1S U31854 ( .A(gray_img[1101]), .B(n28490), .CI(n28489), .CO(n28491) );
  MXL2HS U31855 ( .A(gray_img[1230]), .B(gray_img[1102]), .S(n28507), .OB(
        n28522) );
  INV1S U31856 ( .I(gray_img[1221]), .O(n28502) );
  INV1S U31857 ( .I(gray_img[1220]), .O(n28500) );
  INV1S U31858 ( .I(gray_img[1219]), .O(n28498) );
  INV1S U31859 ( .I(gray_img[1218]), .O(n28496) );
  FA1S U31860 ( .A(gray_img[1089]), .B(gray_img[1088]), .CI(intadd_77_CI), 
        .CO(n28495) );
  FA1S U31861 ( .A(n28496), .B(gray_img[1090]), .CI(n28495), .CO(n28497) );
  FA1S U31862 ( .A(n28498), .B(gray_img[1091]), .CI(n28497), .CO(n28499) );
  FA1S U31863 ( .A(n28500), .B(gray_img[1092]), .CI(n28499), .CO(n28501) );
  MXL2HS U31864 ( .A(gray_img[1229]), .B(gray_img[1101]), .S(n28507), .OB(
        n28565) );
  MXL2HS U31865 ( .A(gray_img[1228]), .B(gray_img[1100]), .S(n28507), .OB(
        n28570) );
  MXL2HS U31866 ( .A(gray_img[1227]), .B(gray_img[1099]), .S(n28507), .OB(
        n28575) );
  MXL2HS U31867 ( .A(gray_img[1226]), .B(gray_img[1098]), .S(n28507), .OB(
        n28580) );
  MXL2HS U31868 ( .A(gray_img[1224]), .B(gray_img[1096]), .S(n28507), .OB(
        n28678) );
  MXL2HS U31869 ( .A(gray_img[1225]), .B(gray_img[1097]), .S(n28507), .OB(
        n28593) );
  OR2 U31870 ( .I1(n29680), .I2(n28516), .O(n28677) );
  INV1S U31871 ( .I(n28516), .O(n28517) );
  INV1S U31872 ( .I(n28672), .O(n28674) );
  OAI112HS U31873 ( .C1(n28522), .C2(n28677), .A1(n28521), .B1(n28520), .O(
        n14031) );
  MUX2S U31874 ( .A(n15889), .B(n28533), .S(gray_img[1356]), .O(n28524) );
  MUX2S U31875 ( .A(n27447), .B(n28533), .S(gray_img[1352]), .O(n28527) );
  AO12S U31876 ( .B1(n15888), .B2(n28536), .A1(n28527), .O(n13993) );
  MUX2S U31877 ( .A(n15889), .B(n28558), .S(gray_img[1484]), .O(n28529) );
  MUX2S U31878 ( .A(n27447), .B(n28558), .S(gray_img[1483]), .O(n28531) );
  ND2S U31879 ( .I1(n15891), .I2(n28581), .O(n28538) );
  OAI112HS U31880 ( .C1(n28585), .C2(n28540), .A1(n28539), .B1(n28538), .O(
        n28541) );
  OAI112HS U31881 ( .C1(n28585), .C2(n28545), .A1(n28544), .B1(n28543), .O(
        n28546) );
  OAI112HS U31882 ( .C1(n28585), .C2(n28550), .A1(n28549), .B1(n28548), .O(
        n28551) );
  OAI112HS U31883 ( .C1(n28585), .C2(n28555), .A1(n28554), .B1(n28553), .O(
        n28556) );
  MUX2S U31884 ( .A(n27447), .B(n28558), .S(gray_img[1480]), .O(n28559) );
  AO12S U31885 ( .B1(n15888), .B2(n28560), .A1(n28559), .O(n13950) );
  OAI112HS U31886 ( .C1(n28565), .C2(n28677), .A1(n28564), .B1(n28563), .O(
        n14032) );
  OAI112HS U31887 ( .C1(n28570), .C2(n28677), .A1(n28569), .B1(n28568), .O(
        n14033) );
  OAI112HS U31888 ( .C1(n28575), .C2(n28677), .A1(n28574), .B1(n28573), .O(
        n14034) );
  OAI112HS U31889 ( .C1(n28580), .C2(n28677), .A1(n28579), .B1(n28578), .O(
        n14035) );
  OAI112HS U31890 ( .C1(n28585), .C2(n28584), .A1(n28583), .B1(n28582), .O(
        n28586) );
  OAI112HS U31891 ( .C1(n28593), .C2(n28677), .A1(n28592), .B1(n28591), .O(
        n14036) );
  MUX2S U31892 ( .A(n15889), .B(n28594), .S(gray_img[1360]), .O(n28595) );
  AO12S U31893 ( .B1(n15888), .B2(n28596), .A1(n28595), .O(n13992) );
  INV1S U31894 ( .I(n28597), .O(n28600) );
  MUX2S U31895 ( .A(gray_img[1360]), .B(gray_img[1488]), .S(n28598), .O(n28599) );
  ND2S U31896 ( .I1(n28600), .I2(n28599), .O(n28604) );
  ND2S U31897 ( .I1(n15888), .I2(n28601), .O(n28602) );
  FA1S U31898 ( .A(intadd_137_B_0_), .B(intadd_137_A_0_), .CI(gray_img[681]), 
        .CO(n28608) );
  FA1S U31899 ( .A(gray_img[682]), .B(n28609), .CI(n28608), .CO(n28610) );
  FA1S U31900 ( .A(gray_img[683]), .B(n28611), .CI(n28610), .CO(n28612) );
  MXL2HS U31901 ( .A(gray_img[558]), .B(gray_img[686]), .S(n28633), .OB(n28648) );
  FA1S U31902 ( .A(gray_img[673]), .B(gray_img[672]), .CI(n28620), .CO(n28621)
         );
  FA1S U31903 ( .A(n28624), .B(gray_img[675]), .CI(n28623), .CO(n28625) );
  MXL2HS U31904 ( .A(gray_img[557]), .B(gray_img[685]), .S(n28633), .OB(n28653) );
  MXL2HS U31905 ( .A(gray_img[556]), .B(gray_img[684]), .S(n28633), .OB(n28658) );
  MXL2HS U31906 ( .A(gray_img[555]), .B(gray_img[683]), .S(n28633), .OB(n28663) );
  MXL2HS U31907 ( .A(gray_img[554]), .B(gray_img[682]), .S(n28633), .OB(n28668) );
  MXL2HS U31908 ( .A(gray_img[552]), .B(gray_img[680]), .S(n28633), .OB(n28684) );
  MXL2HS U31909 ( .A(gray_img[553]), .B(gray_img[681]), .S(n28633), .OB(n28713) );
  INV1S U31910 ( .I(n28642), .O(n28643) );
  OA12S U31911 ( .B1(gray_img[278]), .B2(n29427), .A1(n28707), .O(n28645) );
  MOAI1S U31912 ( .A1(n28707), .A2(gray_img[278]), .B1(n29825), .B2(n28645), 
        .O(n28646) );
  OAI112HS U31913 ( .C1(n28648), .C2(n28712), .A1(n28647), .B1(n28646), .O(
        n13675) );
  ND2S U31914 ( .I1(n28706), .I2(n28649), .O(n28652) );
  INV1S U31915 ( .I(n28707), .O(n28709) );
  OAI112HS U31916 ( .C1(n28653), .C2(n28712), .A1(n28652), .B1(n28651), .O(
        n13676) );
  ND2S U31917 ( .I1(n28706), .I2(n28654), .O(n28657) );
  OAI112HS U31918 ( .C1(n28658), .C2(n28712), .A1(n28657), .B1(n28656), .O(
        n13677) );
  ND2S U31919 ( .I1(n28706), .I2(n28659), .O(n28662) );
  OAI112HS U31920 ( .C1(n28663), .C2(n28712), .A1(n28662), .B1(n28661), .O(
        n13678) );
  ND2S U31921 ( .I1(n28706), .I2(n28664), .O(n28667) );
  OAI112HS U31922 ( .C1(n28668), .C2(n28712), .A1(n28667), .B1(n28666), .O(
        n13679) );
  MUX2S U31923 ( .A(gray_img[1216]), .B(gray_img[1088]), .S(n28669), .O(n28670) );
  OAI112HS U31924 ( .C1(n28678), .C2(n28677), .A1(n28676), .B1(n28675), .O(
        n13742) );
  MUX2S U31925 ( .A(gray_img[544]), .B(gray_img[672]), .S(n28679), .O(n28680)
         );
  ND2S U31926 ( .I1(n28706), .I2(n28680), .O(n28683) );
  OAI112HS U31927 ( .C1(n28684), .C2(n28712), .A1(n28683), .B1(n28682), .O(
        n13784) );
  OA12S U31928 ( .B1(n29831), .B2(n28809), .A1(n28686), .O(n28687) );
  OAI112HS U31929 ( .C1(n28689), .C2(n28812), .A1(n28688), .B1(n28687), .O(
        n15269) );
  OA12S U31930 ( .B1(n29837), .B2(n28809), .A1(n28691), .O(n28692) );
  OAI112HS U31931 ( .C1(n28694), .C2(n28812), .A1(n28693), .B1(n28692), .O(
        n14873) );
  OA12S U31932 ( .B1(n29843), .B2(n28809), .A1(n28696), .O(n28697) );
  OAI112HS U31933 ( .C1(n28699), .C2(n28812), .A1(n28698), .B1(n28697), .O(
        n14673) );
  OA12S U31934 ( .B1(n29849), .B2(n28809), .A1(n28701), .O(n28702) );
  OAI112HS U31935 ( .C1(n28704), .C2(n28812), .A1(n28703), .B1(n28702), .O(
        n14472) );
  ND2S U31936 ( .I1(n28706), .I2(n28705), .O(n28711) );
  OAI112HS U31937 ( .C1(n28713), .C2(n28712), .A1(n28711), .B1(n28710), .O(
        n14469) );
  MUX2S U31938 ( .A(gray_img[2040]), .B(gray_img[1912]), .S(n28715), .O(n28716) );
  ND2S U31939 ( .I1(n28717), .I2(n28716), .O(n28721) );
  ND2S U31940 ( .I1(n15888), .I2(n28718), .O(n28719) );
  ND3S U31941 ( .I1(n28721), .I2(n28720), .I3(n28719), .O(n28722) );
  MUX2S U31942 ( .A(gray_img[952]), .B(gray_img[824]), .S(n28725), .O(n28726)
         );
  OAI112HS U31943 ( .C1(n28734), .C2(n28733), .A1(n28732), .B1(n28731), .O(
        n13775) );
  FA1S U31944 ( .A(gray_img[273]), .B(gray_img[272]), .CI(intadd_169_CI), .CO(
        n28735) );
  FA1S U31945 ( .A(n28736), .B(gray_img[274]), .CI(n28735), .CO(n28737) );
  FA1S U31946 ( .A(n28738), .B(gray_img[275]), .CI(n28737), .CO(n28739) );
  INV1S U31947 ( .I(gray_img[415]), .O(n28764) );
  INV1S U31948 ( .I(gray_img[287]), .O(n28762) );
  INV1S U31949 ( .I(gray_img[412]), .O(n28752) );
  INV1S U31950 ( .I(gray_img[411]), .O(n28750) );
  INV1S U31951 ( .I(gray_img[410]), .O(n28748) );
  FA1S U31952 ( .A(gray_img[281]), .B(gray_img[280]), .CI(intadd_206_CI), .CO(
        n28747) );
  FA1S U31953 ( .A(n28748), .B(gray_img[282]), .CI(n28747), .CO(n28749) );
  INV1S U31954 ( .I(n28756), .O(n28755) );
  INV1S U31955 ( .I(gray_img[285]), .O(n28754) );
  INV1S U31956 ( .I(gray_img[414]), .O(n28753) );
  MOAI1S U31957 ( .A1(n28755), .A2(n28754), .B1(gray_img[286]), .B2(n28753), 
        .O(n28760) );
  NR2 U31958 ( .I1(gray_img[285]), .I2(n28756), .O(n28757) );
  NR2 U31959 ( .I1(gray_img[413]), .I2(n28757), .O(n28759) );
  INV1S U31960 ( .I(gray_img[286]), .O(n28758) );
  MOAI1S U31961 ( .A1(n28760), .A2(n28759), .B1(gray_img[414]), .B2(n28758), 
        .O(n28761) );
  OAI12HS U31962 ( .B1(gray_img[415]), .B2(n28762), .A1(n28761), .O(n28763) );
  OAI12HS U31963 ( .B1(gray_img[287]), .B2(n28764), .A1(n28763), .O(n28765) );
  MXL2HS U31964 ( .A(gray_img[286]), .B(gray_img[414]), .S(n28765), .OB(n28778) );
  MXL2HS U31965 ( .A(gray_img[285]), .B(gray_img[413]), .S(n28765), .OB(n28783) );
  MXL2HS U31966 ( .A(gray_img[284]), .B(gray_img[412]), .S(n28765), .OB(n28788) );
  MXL2HS U31967 ( .A(gray_img[283]), .B(gray_img[411]), .S(n28765), .OB(n28793) );
  MXL2HS U31968 ( .A(gray_img[282]), .B(gray_img[410]), .S(n28765), .OB(n28798) );
  MXL2HS U31969 ( .A(gray_img[280]), .B(gray_img[408]), .S(n28765), .OB(n28817) );
  MXL2HS U31970 ( .A(gray_img[281]), .B(gray_img[409]), .S(n28765), .OB(n28843) );
  INV1S U31971 ( .I(n28775), .O(n28774) );
  NR2 U31972 ( .I1(n29680), .I2(n28774), .O(n28847) );
  OR2 U31973 ( .I1(n29680), .I2(n28775), .O(n28844) );
  MUX2S U31974 ( .A(n15904), .B(n28840), .S(gray_img[142]), .O(n28777) );
  ND2S U31975 ( .I1(n15890), .I2(n28840), .O(n28776) );
  OAI112HS U31976 ( .C1(n28844), .C2(n28778), .A1(n28777), .B1(n28776), .O(
        n28779) );
  OAI112HS U31977 ( .C1(n28844), .C2(n28783), .A1(n28782), .B1(n28781), .O(
        n28784) );
  OAI112HS U31978 ( .C1(n28844), .C2(n28788), .A1(n28787), .B1(n28786), .O(
        n28789) );
  OAI112HS U31979 ( .C1(n28844), .C2(n28793), .A1(n28792), .B1(n28791), .O(
        n28794) );
  OAI112HS U31980 ( .C1(n28844), .C2(n28798), .A1(n28797), .B1(n28796), .O(
        n28799) );
  AO12S U31981 ( .B1(n15888), .B2(n28803), .A1(n28802), .O(n13822) );
  MUX2S U31982 ( .A(gray_img[928]), .B(gray_img[800]), .S(n28804), .O(n28805)
         );
  OA12S U31983 ( .B1(n29734), .B2(n28809), .A1(n28808), .O(n28810) );
  OAI112HS U31984 ( .C1(n28813), .C2(n28812), .A1(n28811), .B1(n28810), .O(
        n13776) );
  MUX2S U31985 ( .A(gray_img[400]), .B(gray_img[272]), .S(n28814), .O(n28819)
         );
  OAI112HS U31986 ( .C1(n28844), .C2(n28817), .A1(n28816), .B1(n28815), .O(
        n28818) );
  ND2S U31987 ( .I1(n26445), .I2(n30081), .O(n28820) );
  OAI112HS U31988 ( .C1(n30077), .C2(n28822), .A1(n28821), .B1(n28820), .O(
        n28823) );
  OAI112HS U31989 ( .C1(n30077), .C2(n28827), .A1(n28826), .B1(n28825), .O(
        n28828) );
  OAI112HS U31990 ( .C1(n30077), .C2(n28832), .A1(n28831), .B1(n28830), .O(
        n28833) );
  OAI112HS U31991 ( .C1(n30077), .C2(n28837), .A1(n28836), .B1(n28835), .O(
        n28838) );
  OAI112HS U31992 ( .C1(n28844), .C2(n28843), .A1(n28842), .B1(n28841), .O(
        n28845) );
  OAI112HS U31993 ( .C1(n30077), .C2(n28850), .A1(n28849), .B1(n28848), .O(
        n28851) );
  INV1S U31994 ( .I(gray_img[1214]), .O(n28863) );
  INV1S U31995 ( .I(gray_img[1213]), .O(n28861) );
  INV1S U31996 ( .I(gray_img[1212]), .O(n28859) );
  INV1S U31997 ( .I(gray_img[1211]), .O(n28857) );
  INV1S U31998 ( .I(gray_img[1210]), .O(n28855) );
  INV1S U31999 ( .I(gray_img[1209]), .O(n28853) );
  INV1S U32000 ( .I(gray_img[1206]), .O(n28876) );
  INV1S U32001 ( .I(gray_img[1205]), .O(n28874) );
  INV1S U32002 ( .I(gray_img[1204]), .O(n28872) );
  INV1S U32003 ( .I(gray_img[1203]), .O(n28870) );
  INV1S U32004 ( .I(gray_img[1202]), .O(n28868) );
  INV1S U32005 ( .I(gray_img[1201]), .O(n28866) );
  FA1S U32006 ( .A(n28868), .B(gray_img[1074]), .CI(n28867), .CO(n28869) );
  MXL2HS U32007 ( .A(gray_img[1206]), .B(gray_img[1078]), .S(n28935), .OB(
        n28892) );
  MXL2HS U32008 ( .A(gray_img[1205]), .B(gray_img[1077]), .S(n28935), .OB(
        n28902) );
  MXL2HS U32009 ( .A(gray_img[1204]), .B(gray_img[1076]), .S(n28935), .OB(
        n28922) );
  MXL2HS U32010 ( .A(gray_img[1203]), .B(gray_img[1075]), .S(n28935), .OB(
        n28927) );
  MXL2HS U32011 ( .A(gray_img[1202]), .B(gray_img[1074]), .S(n28935), .OB(
        n28932) );
  MUX2S U32012 ( .A(gray_img[1209]), .B(gray_img[1081]), .S(n28879), .O(n28949) );
  MXL2HS U32013 ( .A(gray_img[1201]), .B(gray_img[1073]), .S(n28935), .OB(
        n28946) );
  INV1S U32014 ( .I(n28889), .O(n28888) );
  NR2 U32015 ( .I1(n29680), .I2(n28888), .O(n28950) );
  ND2S U32016 ( .I1(n15890), .I2(n28943), .O(n28890) );
  OAI112HS U32017 ( .C1(n28947), .C2(n28892), .A1(n28891), .B1(n28890), .O(
        n28893) );
  ND2S U32018 ( .I1(n27751), .I2(n29344), .O(n28895) );
  OAI112HS U32019 ( .C1(n29340), .C2(n28897), .A1(n28896), .B1(n28895), .O(
        n28898) );
  ND2S U32020 ( .I1(n15891), .I2(n28943), .O(n28900) );
  OAI112HS U32021 ( .C1(n28947), .C2(n28902), .A1(n28901), .B1(n28900), .O(
        n28903) );
  OAI112HS U32022 ( .C1(n29340), .C2(n28907), .A1(n28906), .B1(n28905), .O(
        n28908) );
  OAI112HS U32023 ( .C1(n29340), .C2(n28912), .A1(n28911), .B1(n28910), .O(
        n28913) );
  OAI112HS U32024 ( .C1(n29340), .C2(n28917), .A1(n28916), .B1(n28915), .O(
        n28918) );
  OAI112HS U32025 ( .C1(n28947), .C2(n28922), .A1(n28921), .B1(n28920), .O(
        n28923) );
  OAI112HS U32026 ( .C1(n28947), .C2(n28927), .A1(n28926), .B1(n28925), .O(
        n28928) );
  OAI112HS U32027 ( .C1(n28947), .C2(n28932), .A1(n28931), .B1(n28930), .O(
        n28933) );
  INV1S U32028 ( .I(n28947), .O(n28937) );
  MUX2S U32029 ( .A(gray_img[1200]), .B(gray_img[1072]), .S(n28935), .O(n28936) );
  ND2S U32030 ( .I1(n28937), .I2(n28936), .O(n28940) );
  MUX2S U32031 ( .A(n29032), .B(n28943), .S(gray_img[536]), .O(n28939) );
  ND2S U32032 ( .I1(n15888), .I2(n28943), .O(n28938) );
  OAI112HS U32033 ( .C1(n28947), .C2(n28946), .A1(n28945), .B1(n28944), .O(
        n28948) );
  INV1S U32034 ( .I(gray_img[1447]), .O(n28962) );
  INV1S U32035 ( .I(gray_img[1445]), .O(n28958) );
  INV1S U32036 ( .I(gray_img[1444]), .O(n28956) );
  INV1S U32037 ( .I(gray_img[1443]), .O(n28954) );
  FA1S U32038 ( .A(gray_img[1313]), .B(gray_img[1312]), .CI(intadd_60_CI), 
        .CO(n28951) );
  FA1S U32039 ( .A(n28952), .B(gray_img[1314]), .CI(n28951), .CO(n28953) );
  FA1S U32040 ( .A(n28954), .B(gray_img[1315]), .CI(n28953), .CO(n28955) );
  FA1S U32041 ( .A(n28956), .B(gray_img[1316]), .CI(n28955), .CO(n28957) );
  MXL2HS U32042 ( .A(gray_img[1446]), .B(gray_img[1318]), .S(n29009), .OB(
        n28986) );
  INV1S U32043 ( .I(gray_img[1454]), .O(n28972) );
  INV1S U32044 ( .I(gray_img[1452]), .O(n28968) );
  INV1S U32045 ( .I(gray_img[1450]), .O(n28964) );
  FA1S U32046 ( .A(gray_img[1321]), .B(gray_img[1320]), .CI(intadd_59_CI), 
        .CO(n28963) );
  MXL2HS U32047 ( .A(gray_img[1445]), .B(gray_img[1317]), .S(n29009), .OB(
        n28991) );
  MXL2HS U32048 ( .A(gray_img[1444]), .B(gray_img[1316]), .S(n29009), .OB(
        n28996) );
  MXL2HS U32049 ( .A(gray_img[1443]), .B(gray_img[1315]), .S(n29009), .OB(
        n29001) );
  MXL2HS U32050 ( .A(gray_img[1442]), .B(gray_img[1314]), .S(n29009), .OB(
        n29006) );
  MXL2HS U32051 ( .A(gray_img[1441]), .B(gray_img[1313]), .S(n29009), .OB(
        n29036) );
  FA1S U32052 ( .A(n29016), .B(n29036), .CI(n29039), .CO(n28976) );
  INV1S U32053 ( .I(n28983), .O(n28982) );
  NR2 U32054 ( .I1(n29680), .I2(n28982), .O(n29040) );
  OR2 U32055 ( .I1(n29680), .I2(n28983), .O(n29037) );
  ND2S U32056 ( .I1(n15890), .I2(n29033), .O(n28984) );
  OAI112HS U32057 ( .C1(n29037), .C2(n28986), .A1(n28985), .B1(n28984), .O(
        n28987) );
  OAI112HS U32058 ( .C1(n29037), .C2(n28991), .A1(n28990), .B1(n28989), .O(
        n28992) );
  OAI112HS U32059 ( .C1(n29037), .C2(n28996), .A1(n28995), .B1(n28994), .O(
        n28997) );
  OAI112HS U32060 ( .C1(n29037), .C2(n29001), .A1(n29000), .B1(n28999), .O(
        n29002) );
  OAI112HS U32061 ( .C1(n29037), .C2(n29006), .A1(n29005), .B1(n29004), .O(
        n29007) );
  INV1S U32062 ( .I(n29037), .O(n29011) );
  MUX2S U32063 ( .A(gray_img[1440]), .B(gray_img[1312]), .S(n29009), .O(n29010) );
  ND2S U32064 ( .I1(n29011), .I2(n29010), .O(n29014) );
  MUX2S U32065 ( .A(n30005), .B(n29033), .S(gray_img[656]), .O(n29013) );
  ND2S U32066 ( .I1(n15888), .I2(n29033), .O(n29012) );
  ND3S U32067 ( .I1(n29014), .I2(n29013), .I3(n29012), .O(n29015) );
  OA12S U32068 ( .B1(n29831), .B2(n29046), .A1(n29018), .O(n29019) );
  OAI112HS U32069 ( .C1(n29021), .C2(n29049), .A1(n29020), .B1(n29019), .O(
        n14050) );
  OA12S U32070 ( .B1(n29837), .B2(n29046), .A1(n29023), .O(n29024) );
  OAI112HS U32071 ( .C1(n29026), .C2(n29049), .A1(n29025), .B1(n29024), .O(
        n14051) );
  OA12S U32072 ( .B1(n29843), .B2(n29046), .A1(n29028), .O(n29029) );
  OAI112HS U32073 ( .C1(n29031), .C2(n29049), .A1(n29030), .B1(n29029), .O(
        n14052) );
  OAI112HS U32074 ( .C1(n29037), .C2(n29036), .A1(n29035), .B1(n29034), .O(
        n29038) );
  MUX2S U32075 ( .A(gray_img[1192]), .B(gray_img[1064]), .S(n29041), .O(n29042) );
  OA12S U32076 ( .B1(n29734), .B2(n29046), .A1(n29045), .O(n29047) );
  OAI112HS U32077 ( .C1(n29050), .C2(n29049), .A1(n29048), .B1(n29047), .O(
        n13744) );
  MAO222S U32078 ( .A1(gray_img[657]), .B1(gray_img[656]), .C1(n29051), .O(
        n29052) );
  INV1S U32079 ( .I(gray_img[540]), .O(n29070) );
  INV1S U32080 ( .I(gray_img[538]), .O(n29066) );
  FA1S U32081 ( .A(n29064), .B(gray_img[665]), .CI(n29063), .CO(n29065) );
  ND2S U32082 ( .I1(n29071), .I2(gray_img[541]), .O(n29074) );
  INV1S U32083 ( .I(gray_img[670]), .O(n29072) );
  OAI22S U32084 ( .A1(gray_img[542]), .A2(n29072), .B1(n29071), .B2(
        gray_img[541]), .O(n29073) );
  AOI12HS U32085 ( .B1(n29075), .B2(n29074), .A1(n29073), .O(n29078) );
  NR2 U32086 ( .I1(gray_img[670]), .I2(n29076), .O(n29077) );
  MOAI1S U32087 ( .A1(n29078), .A2(n29077), .B1(gray_img[671]), .B2(n29080), 
        .O(n29079) );
  OAI12HS U32088 ( .B1(gray_img[671]), .B2(n29080), .A1(n29079), .O(n29351) );
  MXL2HS U32089 ( .A(gray_img[670]), .B(gray_img[542]), .S(n29351), .OB(n29094) );
  MXL2HS U32090 ( .A(gray_img[669]), .B(gray_img[541]), .S(n29351), .OB(n29317) );
  MXL2HS U32091 ( .A(gray_img[668]), .B(gray_img[540]), .S(n29351), .OB(n29327) );
  MXL2HS U32092 ( .A(gray_img[667]), .B(gray_img[539]), .S(n29351), .OB(n29332) );
  MXL2HS U32093 ( .A(gray_img[666]), .B(gray_img[538]), .S(n29351), .OB(n29337) );
  MXL2HS U32094 ( .A(gray_img[665]), .B(gray_img[537]), .S(n29351), .OB(n29377) );
  INV1S U32095 ( .I(n29091), .O(n29090) );
  NR2 U32096 ( .I1(n29680), .I2(n29090), .O(n29381) );
  OR2 U32097 ( .I1(n29680), .I2(n29091), .O(n29378) );
  ND2S U32098 ( .I1(n15890), .I2(n29374), .O(n29092) );
  OAI112HS U32099 ( .C1(n29378), .C2(n29094), .A1(n29093), .B1(n29092), .O(
        n29095) );
  INV1S U32100 ( .I(gray_img[1709]), .O(n29104) );
  INV1S U32101 ( .I(gray_img[1707]), .O(n29100) );
  INV1S U32102 ( .I(gray_img[1706]), .O(n29098) );
  FA1S U32103 ( .A(gray_img[1577]), .B(gray_img[1576]), .CI(intadd_47_CI), 
        .CO(n29097) );
  FA1S U32104 ( .A(n29098), .B(gray_img[1578]), .CI(n29097), .CO(n29099) );
  FA1S U32105 ( .A(n29100), .B(gray_img[1579]), .CI(n29099), .CO(n29101) );
  FA1S U32106 ( .A(n29102), .B(gray_img[1580]), .CI(n29101), .CO(n29103) );
  INV1S U32107 ( .I(gray_img[1703]), .O(n29120) );
  INV1S U32108 ( .I(gray_img[1702]), .O(n29118) );
  INV1S U32109 ( .I(gray_img[1701]), .O(n29116) );
  INV1S U32110 ( .I(gray_img[1700]), .O(n29114) );
  INV1S U32111 ( .I(gray_img[1699]), .O(n29112) );
  INV1S U32112 ( .I(gray_img[1698]), .O(n29110) );
  MAO222S U32113 ( .A1(gray_img[1569]), .B1(gray_img[1568]), .C1(intadd_48_CI), 
        .O(n29109) );
  FA1S U32114 ( .A(n29110), .B(gray_img[1570]), .CI(n29109), .CO(n29111) );
  FA1S U32115 ( .A(n29112), .B(gray_img[1571]), .CI(n29111), .CO(n29113) );
  FA1S U32116 ( .A(n29114), .B(gray_img[1572]), .CI(n29113), .CO(n29115) );
  FA1S U32117 ( .A(n29116), .B(gray_img[1573]), .CI(n29115), .CO(n29117) );
  MXL2HS U32118 ( .A(gray_img[1702]), .B(gray_img[1574]), .S(n29183), .OB(
        n29134) );
  MXL2HS U32119 ( .A(gray_img[1701]), .B(gray_img[1573]), .S(n29183), .OB(
        n29139) );
  MXL2HS U32120 ( .A(gray_img[1700]), .B(gray_img[1572]), .S(n29183), .OB(
        n29144) );
  MXL2HS U32121 ( .A(gray_img[1699]), .B(gray_img[1571]), .S(n29183), .OB(
        n29149) );
  MXL2HS U32122 ( .A(gray_img[1698]), .B(gray_img[1570]), .S(n29183), .OB(
        n29154) );
  MXL2HS U32123 ( .A(gray_img[1697]), .B(gray_img[1569]), .S(n29183), .OB(
        n29159) );
  INV1S U32124 ( .I(n29131), .O(n29130) );
  NR2 U32125 ( .I1(n29680), .I2(n29130), .O(n29192) );
  OR2 U32126 ( .I1(n29680), .I2(n29131), .O(n29182) );
  MUX2S U32127 ( .A(n29587), .B(n29186), .S(gray_img[790]), .O(n29133) );
  ND2S U32128 ( .I1(n15890), .I2(n29186), .O(n29132) );
  OAI112HS U32129 ( .C1(n29182), .C2(n29134), .A1(n29133), .B1(n29132), .O(
        n29135) );
  MUX2S U32130 ( .A(n15904), .B(n29186), .S(gray_img[789]), .O(n29138) );
  OAI112HS U32131 ( .C1(n29182), .C2(n29139), .A1(n29138), .B1(n29137), .O(
        n29140) );
  OAI112HS U32132 ( .C1(n29182), .C2(n29144), .A1(n29143), .B1(n29142), .O(
        n29145) );
  OAI112HS U32133 ( .C1(n29182), .C2(n29149), .A1(n29148), .B1(n29147), .O(
        n29150) );
  OAI112HS U32134 ( .C1(n29182), .C2(n29154), .A1(n29153), .B1(n29152), .O(
        n29155) );
  OAI112HS U32135 ( .C1(n29182), .C2(n29159), .A1(n29158), .B1(n29157), .O(
        n29160) );
  INV1S U32136 ( .I(n30021), .O(n30023) );
  OAI112HS U32137 ( .C1(n29166), .C2(n30026), .A1(n29165), .B1(n29164), .O(
        n13830) );
  OAI112HS U32138 ( .C1(n29171), .C2(n30026), .A1(n29170), .B1(n29169), .O(
        n13630) );
  OAI112HS U32139 ( .C1(n29176), .C2(n30026), .A1(n29175), .B1(n29174), .O(
        n13640) );
  OAI112HS U32140 ( .C1(n29181), .C2(n30026), .A1(n29180), .B1(n29179), .O(
        n13661) );
  INV1S U32141 ( .I(n29182), .O(n29185) );
  MUX2S U32142 ( .A(gray_img[1696]), .B(gray_img[1568]), .S(n29183), .O(n29184) );
  ND2S U32143 ( .I1(n29185), .I2(n29184), .O(n29189) );
  ND2S U32144 ( .I1(n15888), .I2(n29186), .O(n29187) );
  ND3S U32145 ( .I1(n29189), .I2(n29188), .I3(n29187), .O(n29190) );
  OAI112HS U32146 ( .C1(n29197), .C2(n30026), .A1(n29196), .B1(n29195), .O(
        n13685) );
  INV1S U32147 ( .I(gray_img[1726]), .O(n29207) );
  INV1S U32148 ( .I(gray_img[1723]), .O(n29201) );
  INV1S U32149 ( .I(gray_img[1722]), .O(n29199) );
  MAO222S U32150 ( .A1(gray_img[1593]), .B1(gray_img[1592]), .C1(intadd_45_CI), 
        .O(n29198) );
  FA1S U32151 ( .A(n29199), .B(gray_img[1594]), .CI(n29198), .CO(n29200) );
  FA1S U32152 ( .A(n29201), .B(gray_img[1595]), .CI(n29200), .CO(n29202) );
  FA1S U32153 ( .A(n29203), .B(gray_img[1596]), .CI(n29202), .CO(n29204) );
  MXL2HS U32154 ( .A(gray_img[1726]), .B(gray_img[1598]), .S(n29258), .OB(
        n29237) );
  INV1S U32155 ( .I(gray_img[1717]), .O(n29217) );
  INV1S U32156 ( .I(gray_img[1716]), .O(n29215) );
  FA1S U32157 ( .A(gray_img[1585]), .B(gray_img[1584]), .CI(intadd_44_CI), 
        .CO(n29210) );
  FA1S U32158 ( .A(n29211), .B(gray_img[1586]), .CI(n29210), .CO(n29212) );
  FA1S U32159 ( .A(n29213), .B(gray_img[1587]), .CI(n29212), .CO(n29214) );
  FA1S U32160 ( .A(n29215), .B(gray_img[1588]), .CI(n29214), .CO(n29216) );
  MXL2HS U32161 ( .A(gray_img[1725]), .B(gray_img[1597]), .S(n29258), .OB(
        n29240) );
  MXL2HS U32162 ( .A(gray_img[1724]), .B(gray_img[1596]), .S(n29258), .OB(
        n29245) );
  MXL2HS U32163 ( .A(gray_img[1723]), .B(gray_img[1595]), .S(n29258), .OB(
        n29250) );
  MXL2HS U32164 ( .A(gray_img[1722]), .B(gray_img[1594]), .S(n29258), .OB(
        n29255) );
  MXL2HS U32165 ( .A(gray_img[1721]), .B(gray_img[1593]), .S(n29258), .OB(
        n29269) );
  OR2 U32166 ( .I1(n29680), .I2(n29231), .O(n29270) );
  INV1S U32167 ( .I(n29231), .O(n29232) );
  OA12S U32168 ( .B1(gray_img[798]), .B2(n29427), .A1(n29266), .O(n29234) );
  MOAI1S U32169 ( .A1(gray_img[798]), .A2(n29266), .B1(n29825), .B2(n29234), 
        .O(n29235) );
  OAI112HS U32170 ( .C1(n29237), .C2(n29270), .A1(n29236), .B1(n29235), .O(
        n13885) );
  ND2S U32171 ( .I1(n26828), .I2(n29266), .O(n29238) );
  OAI112HS U32172 ( .C1(n29270), .C2(n29240), .A1(n29239), .B1(n29238), .O(
        n29241) );
  OAI112HS U32173 ( .C1(n29270), .C2(n29245), .A1(n29244), .B1(n29243), .O(
        n29246) );
  OAI112HS U32174 ( .C1(n29270), .C2(n29250), .A1(n29249), .B1(n29248), .O(
        n29251) );
  OAI112HS U32175 ( .C1(n29270), .C2(n29255), .A1(n29254), .B1(n29253), .O(
        n29256) );
  INV1S U32176 ( .I(n29270), .O(n29260) );
  MUX2S U32177 ( .A(gray_img[1720]), .B(gray_img[1592]), .S(n29258), .O(n29259) );
  ND2S U32178 ( .I1(n29260), .I2(n29259), .O(n29263) );
  ND2S U32179 ( .I1(n15888), .I2(n29266), .O(n29261) );
  ND3S U32180 ( .I1(n29263), .I2(n29262), .I3(n29261), .O(n29264) );
  OAI112HS U32181 ( .C1(n29270), .C2(n29269), .A1(n29268), .B1(n29267), .O(
        n29271) );
  INV1S U32182 ( .I(gray_img[926]), .O(n29284) );
  INV1S U32183 ( .I(gray_img[924]), .O(n29280) );
  INV1S U32184 ( .I(gray_img[923]), .O(n29278) );
  INV1S U32185 ( .I(gray_img[919]), .O(n29298) );
  INV1S U32186 ( .I(gray_img[918]), .O(n29296) );
  INV1S U32187 ( .I(gray_img[917]), .O(n29294) );
  INV1S U32188 ( .I(gray_img[916]), .O(n29292) );
  INV1S U32189 ( .I(gray_img[915]), .O(n29290) );
  INV1S U32190 ( .I(gray_img[914]), .O(n29288) );
  FA1S U32191 ( .A(gray_img[784]), .B(gray_img[785]), .CI(intadd_156_CI), .CO(
        n29287) );
  FA1S U32192 ( .A(n29288), .B(gray_img[786]), .CI(n29287), .CO(n29289) );
  FA1S U32193 ( .A(n29290), .B(gray_img[787]), .CI(n29289), .CO(n29291) );
  FA1S U32194 ( .A(n29292), .B(gray_img[788]), .CI(n29291), .CO(n29293) );
  FA1S U32195 ( .A(n29294), .B(gray_img[789]), .CI(n29293), .CO(n29295) );
  MXL2HS U32196 ( .A(gray_img[918]), .B(gray_img[790]), .S(n30029), .OB(n29312) );
  MXL2HS U32197 ( .A(gray_img[917]), .B(gray_img[789]), .S(n30029), .OB(n29322) );
  MXL2HS U32198 ( .A(gray_img[916]), .B(gray_img[788]), .S(n30029), .OB(n29361) );
  MXL2HS U32199 ( .A(gray_img[915]), .B(gray_img[787]), .S(n30029), .OB(n29366) );
  MXL2HS U32200 ( .A(gray_img[914]), .B(gray_img[786]), .S(n30029), .OB(n29371) );
  MUX2S U32201 ( .A(gray_img[920]), .B(gray_img[792]), .S(n29299), .O(n30037)
         );
  MXL2HS U32202 ( .A(gray_img[913]), .B(gray_img[785]), .S(n30029), .OB(n29384) );
  MUX2S U32203 ( .A(gray_img[921]), .B(gray_img[793]), .S(n29299), .O(n29386)
         );
  INV1S U32204 ( .I(n29309), .O(n29308) );
  NR2 U32205 ( .I1(n29680), .I2(n29308), .O(n30038) );
  OR2 U32206 ( .I1(n29680), .I2(n29309), .O(n30028) );
  ND2S U32207 ( .I1(n15890), .I2(n30032), .O(n29310) );
  OAI112HS U32208 ( .C1(n30028), .C2(n29312), .A1(n29311), .B1(n29310), .O(
        n29313) );
  ND2S U32209 ( .I1(n26445), .I2(n29374), .O(n29315) );
  OAI112HS U32210 ( .C1(n29378), .C2(n29317), .A1(n29316), .B1(n29315), .O(
        n29318) );
  ND2S U32211 ( .I1(n15891), .I2(n30032), .O(n29320) );
  OAI112HS U32212 ( .C1(n30028), .C2(n29322), .A1(n29321), .B1(n29320), .O(
        n29323) );
  OAI112HS U32213 ( .C1(n29378), .C2(n29327), .A1(n29326), .B1(n29325), .O(
        n29328) );
  OAI112HS U32214 ( .C1(n29378), .C2(n29332), .A1(n29331), .B1(n29330), .O(
        n29333) );
  OAI112HS U32215 ( .C1(n29378), .C2(n29337), .A1(n29336), .B1(n29335), .O(
        n29338) );
  INV1S U32216 ( .I(n29340), .O(n29343) );
  MUX2S U32217 ( .A(gray_img[1464]), .B(gray_img[1336]), .S(n29341), .O(n29342) );
  ND2S U32218 ( .I1(n29343), .I2(n29342), .O(n29347) );
  ND2S U32219 ( .I1(n15888), .I2(n29344), .O(n29345) );
  ND3S U32220 ( .I1(n29347), .I2(n29346), .I3(n29345), .O(n29348) );
  INV1S U32221 ( .I(n29378), .O(n29353) );
  MUX2S U32222 ( .A(gray_img[664]), .B(gray_img[536]), .S(n29351), .O(n29352)
         );
  ND2S U32223 ( .I1(n29353), .I2(n29352), .O(n29356) );
  ND2S U32224 ( .I1(n15888), .I2(n29374), .O(n29354) );
  ND3S U32225 ( .I1(n29356), .I2(n29355), .I3(n29354), .O(n29357) );
  OAI112HS U32226 ( .C1(n30028), .C2(n29361), .A1(n29360), .B1(n29359), .O(
        n29362) );
  OAI112HS U32227 ( .C1(n30028), .C2(n29366), .A1(n29365), .B1(n29364), .O(
        n29367) );
  OAI112HS U32228 ( .C1(n30028), .C2(n29371), .A1(n29370), .B1(n29369), .O(
        n29372) );
  OAI112HS U32229 ( .C1(n29378), .C2(n29377), .A1(n29376), .B1(n29375), .O(
        n29379) );
  OAI112HS U32230 ( .C1(n30028), .C2(n29384), .A1(n29383), .B1(n29382), .O(
        n29385) );
  INV1S U32231 ( .I(gray_img[1796]), .O(n29393) );
  INV1S U32232 ( .I(gray_img[1795]), .O(n29391) );
  INV1S U32233 ( .I(gray_img[1793]), .O(n29387) );
  MXL2HS U32234 ( .A(gray_img[1798]), .B(gray_img[1926]), .S(n30089), .OB(
        n29431) );
  FA1S U32235 ( .A(gray_img[1800]), .B(n29400), .CI(gray_img[1801]), .CO(
        n29401) );
  ND2S U32236 ( .I1(n29411), .I2(gray_img[1807]), .O(n29412) );
  AOI22S U32237 ( .A1(gray_img[1935]), .A2(n29414), .B1(n29413), .B2(n29412), 
        .O(n29415) );
  MXL2HS U32238 ( .A(gray_img[1797]), .B(gray_img[1925]), .S(n30089), .OB(
        n29459) );
  MXL2HS U32239 ( .A(gray_img[1796]), .B(gray_img[1924]), .S(n30089), .OB(
        n29464) );
  MXL2HS U32240 ( .A(gray_img[1795]), .B(gray_img[1923]), .S(n30089), .OB(
        n29469) );
  MXL2HS U32241 ( .A(gray_img[1794]), .B(gray_img[1922]), .S(n30089), .OB(
        n29474) );
  MXL2HS U32242 ( .A(gray_img[1793]), .B(gray_img[1921]), .S(n30089), .OB(
        n29490) );
  OR2 U32243 ( .I1(n29680), .I2(n29424), .O(n30088) );
  INV1S U32244 ( .I(n29424), .O(n29425) );
  OA12S U32245 ( .B1(gray_img[902]), .B2(n29427), .A1(n30092), .O(n29428) );
  MOAI1S U32246 ( .A1(gray_img[902]), .A2(n30092), .B1(n29825), .B2(n29428), 
        .O(n29429) );
  OAI112HS U32247 ( .C1(n29431), .C2(n30088), .A1(n29430), .B1(n29429), .O(
        n13839) );
  ND2S U32248 ( .I1(n27751), .I2(n29481), .O(n29432) );
  OAI112HS U32249 ( .C1(n29477), .C2(n29434), .A1(n29433), .B1(n29432), .O(
        n29435) );
  OAI112HS U32250 ( .C1(n29477), .C2(n29439), .A1(n29438), .B1(n29437), .O(
        n29440) );
  ND2S U32251 ( .I1(n15887), .I2(n29481), .O(n29442) );
  OAI112HS U32252 ( .C1(n29477), .C2(n29444), .A1(n29443), .B1(n29442), .O(
        n29445) );
  ND2S U32253 ( .I1(n15934), .I2(n29481), .O(n29447) );
  OAI112HS U32254 ( .C1(n29477), .C2(n29449), .A1(n29448), .B1(n29447), .O(
        n29450) );
  ND2S U32255 ( .I1(n15928), .I2(n29481), .O(n29452) );
  OAI112HS U32256 ( .C1(n29477), .C2(n29454), .A1(n29453), .B1(n29452), .O(
        n29455) );
  ND2S U32257 ( .I1(n26828), .I2(n30092), .O(n29457) );
  OAI112HS U32258 ( .C1(n30088), .C2(n29459), .A1(n29458), .B1(n29457), .O(
        n29460) );
  OAI112HS U32259 ( .C1(n30088), .C2(n29464), .A1(n29463), .B1(n29462), .O(
        n29465) );
  OAI112HS U32260 ( .C1(n30088), .C2(n29469), .A1(n29468), .B1(n29467), .O(
        n29470) );
  OAI112HS U32261 ( .C1(n30088), .C2(n29474), .A1(n29473), .B1(n29472), .O(
        n29475) );
  INV1S U32262 ( .I(n29477), .O(n29480) );
  MUX2S U32263 ( .A(gray_img[1536]), .B(gray_img[1664]), .S(n29478), .O(n29479) );
  ND2S U32264 ( .I1(n29480), .I2(n29479), .O(n29484) );
  ND2S U32265 ( .I1(n15888), .I2(n29481), .O(n29482) );
  OAI112HS U32266 ( .C1(n30088), .C2(n29490), .A1(n29489), .B1(n29488), .O(
        n29491) );
  INV1S U32267 ( .I(gray_img[1943]), .O(n29504) );
  INV1S U32268 ( .I(gray_img[1942]), .O(n29502) );
  INV1S U32269 ( .I(gray_img[1941]), .O(n29500) );
  INV1S U32270 ( .I(gray_img[1940]), .O(n29498) );
  INV1S U32271 ( .I(gray_img[1939]), .O(n29496) );
  INV1S U32272 ( .I(gray_img[1938]), .O(n29494) );
  FA1S U32273 ( .A(gray_img[1808]), .B(gray_img[1809]), .CI(intadd_151_CI), 
        .CO(n29493) );
  FA1S U32274 ( .A(n29494), .B(gray_img[1810]), .CI(n29493), .CO(n29495) );
  FA1S U32275 ( .A(n29496), .B(gray_img[1811]), .CI(n29495), .CO(n29497) );
  FA1S U32276 ( .A(n29498), .B(gray_img[1812]), .CI(n29497), .CO(n29499) );
  FA1S U32277 ( .A(n29500), .B(gray_img[1813]), .CI(n29499), .CO(n29501) );
  MXL2HS U32278 ( .A(gray_img[1942]), .B(gray_img[1814]), .S(n29594), .OB(
        n29528) );
  INV1S U32279 ( .I(gray_img[1949]), .O(n29512) );
  INV1S U32280 ( .I(gray_img[1948]), .O(n29510) );
  INV1S U32281 ( .I(gray_img[1946]), .O(n29506) );
  FA1S U32282 ( .A(gray_img[1816]), .B(gray_img[1817]), .CI(intadd_150_CI), 
        .CO(n29505) );
  MXL2HS U32283 ( .A(gray_img[1941]), .B(gray_img[1813]), .S(n29594), .OB(
        n29558) );
  MXL2HS U32284 ( .A(gray_img[1940]), .B(gray_img[1812]), .S(n29594), .OB(
        n29563) );
  MXL2HS U32285 ( .A(gray_img[1939]), .B(gray_img[1811]), .S(n29594), .OB(
        n29569) );
  MXL2HS U32286 ( .A(gray_img[1938]), .B(gray_img[1810]), .S(n29594), .OB(
        n29574) );
  MUX2S U32287 ( .A(gray_img[1945]), .B(gray_img[1817]), .S(n29517), .O(n29592) );
  MXL2HS U32288 ( .A(gray_img[1937]), .B(gray_img[1809]), .S(n29594), .OB(
        n29590) );
  MUX2S U32289 ( .A(gray_img[1944]), .B(gray_img[1816]), .S(n29517), .O(n29603) );
  FA1S U32290 ( .A(n29592), .B(n29590), .CI(n29603), .CO(n29518) );
  INV1S U32291 ( .I(n29525), .O(n29524) );
  NR2 U32292 ( .I1(n29680), .I2(n29524), .O(n29604) );
  OR2 U32293 ( .I1(n29680), .I2(n29525), .O(n29593) );
  ND2S U32294 ( .I1(n15890), .I2(n29598), .O(n29526) );
  OAI112HS U32295 ( .C1(n29593), .C2(n29528), .A1(n29527), .B1(n29526), .O(
        n29529) );
  ND2S U32296 ( .I1(n29579), .I2(n29531), .O(n29534) );
  INV1S U32297 ( .I(n29580), .O(n29582) );
  MUX2S U32298 ( .A(n29597), .B(n29580), .S(gray_img[781]), .O(n29532) );
  OA12S U32299 ( .B1(n29831), .B2(n29582), .A1(n29532), .O(n29533) );
  OAI112HS U32300 ( .C1(n29535), .C2(n29585), .A1(n29534), .B1(n29533), .O(
        n13898) );
  ND2S U32301 ( .I1(n29579), .I2(n29536), .O(n29539) );
  MUX2S U32302 ( .A(n30050), .B(n29580), .S(gray_img[780]), .O(n29537) );
  OA12S U32303 ( .B1(n29837), .B2(n29582), .A1(n29537), .O(n29538) );
  OAI112HS U32304 ( .C1(n29540), .C2(n29585), .A1(n29539), .B1(n29538), .O(
        n13899) );
  ND2S U32305 ( .I1(n29579), .I2(n29541), .O(n29544) );
  MUX2S U32306 ( .A(n29587), .B(n29580), .S(gray_img[779]), .O(n29542) );
  OA12S U32307 ( .B1(n29843), .B2(n29582), .A1(n29542), .O(n29543) );
  OAI112HS U32308 ( .C1(n29545), .C2(n29585), .A1(n29544), .B1(n29543), .O(
        n13649) );
  ND2S U32309 ( .I1(n29579), .I2(n29546), .O(n29549) );
  MUX2S U32310 ( .A(n29566), .B(n29580), .S(gray_img[778]), .O(n29547) );
  OA12S U32311 ( .B1(n29849), .B2(n29582), .A1(n29547), .O(n29548) );
  OAI112HS U32312 ( .C1(n29550), .C2(n29585), .A1(n29549), .B1(n29548), .O(
        n13670) );
  ND2S U32313 ( .I1(n29579), .I2(n29551), .O(n29554) );
  MUX2S U32314 ( .A(n30044), .B(n29580), .S(gray_img[777]), .O(n29552) );
  OA12S U32315 ( .B1(n29884), .B2(n29582), .A1(n29552), .O(n29553) );
  OAI112HS U32316 ( .C1(n29555), .C2(n29585), .A1(n29554), .B1(n29553), .O(
        n13694) );
  OAI112HS U32317 ( .C1(n29593), .C2(n29558), .A1(n29557), .B1(n29556), .O(
        n29559) );
  OAI112HS U32318 ( .C1(n29593), .C2(n29563), .A1(n29562), .B1(n29561), .O(
        n29564) );
  OAI112HS U32319 ( .C1(n29593), .C2(n29569), .A1(n29568), .B1(n29567), .O(
        n29570) );
  OAI112HS U32320 ( .C1(n29593), .C2(n29574), .A1(n29573), .B1(n29572), .O(
        n29575) );
  MUX2S U32321 ( .A(gray_img[1680]), .B(gray_img[1552]), .S(n29577), .O(n29578) );
  ND2S U32322 ( .I1(n29579), .I2(n29578), .O(n29584) );
  MUX2S U32323 ( .A(n29597), .B(n29580), .S(gray_img[776]), .O(n29581) );
  OA12S U32324 ( .B1(n29734), .B2(n29582), .A1(n29581), .O(n29583) );
  OAI112HS U32325 ( .C1(n29586), .C2(n29585), .A1(n29584), .B1(n29583), .O(
        n13721) );
  OAI112HS U32326 ( .C1(n29593), .C2(n29590), .A1(n29589), .B1(n29588), .O(
        n29591) );
  MUX2S U32327 ( .A(gray_img[1936]), .B(gray_img[1808]), .S(n29594), .O(n29595) );
  ND2S U32328 ( .I1(n29596), .I2(n29595), .O(n29601) );
  ND2S U32329 ( .I1(n15888), .I2(n29598), .O(n29599) );
  ND3S U32330 ( .I1(n29601), .I2(n29600), .I3(n29599), .O(n29602) );
  FA1S U32331 ( .A(gray_img[776]), .B(gray_img[777]), .CI(intadd_147_CI), .CO(
        n29605) );
  FA1S U32332 ( .A(n29606), .B(gray_img[778]), .CI(n29605), .CO(n29607) );
  FA1S U32333 ( .A(n29608), .B(gray_img[779]), .CI(n29607), .CO(n29609) );
  INV1S U32334 ( .I(gray_img[902]), .O(n29626) );
  INV1S U32335 ( .I(gray_img[901]), .O(n29624) );
  INV1S U32336 ( .I(gray_img[900]), .O(n29622) );
  INV1S U32337 ( .I(gray_img[899]), .O(n29620) );
  INV1S U32338 ( .I(gray_img[898]), .O(n29618) );
  MXL2HS U32339 ( .A(gray_img[902]), .B(gray_img[774]), .S(n30100), .OB(n29642) );
  MXL2HS U32340 ( .A(gray_img[901]), .B(gray_img[773]), .S(n30100), .OB(n29973) );
  MXL2HS U32341 ( .A(gray_img[900]), .B(gray_img[772]), .S(n30100), .OB(n29978) );
  MXL2HS U32342 ( .A(gray_img[899]), .B(gray_img[771]), .S(n30100), .OB(n29983) );
  MXL2HS U32343 ( .A(gray_img[898]), .B(gray_img[770]), .S(n30100), .OB(n29988) );
  MXL2HS U32344 ( .A(gray_img[897]), .B(gray_img[769]), .S(n30100), .OB(n30015) );
  INV1S U32345 ( .I(n29639), .O(n29638) );
  NR2 U32346 ( .I1(n29680), .I2(n29638), .O(n30109) );
  ND2S U32347 ( .I1(n15890), .I2(n30103), .O(n29640) );
  OAI112HS U32348 ( .C1(n30099), .C2(n29642), .A1(n29641), .B1(n29640), .O(
        n29643) );
  INV1S U32349 ( .I(gray_img[1415]), .O(n29656) );
  INV1S U32350 ( .I(gray_img[1413]), .O(n29652) );
  INV1S U32351 ( .I(gray_img[1411]), .O(n29648) );
  FA1S U32352 ( .A(gray_img[1281]), .B(gray_img[1280]), .CI(intadd_66_CI), 
        .CO(n29645) );
  FA1S U32353 ( .A(n29646), .B(gray_img[1282]), .CI(n29645), .CO(n29647) );
  FA1S U32354 ( .A(n29648), .B(gray_img[1283]), .CI(n29647), .CO(n29649) );
  FA1S U32355 ( .A(n29650), .B(gray_img[1284]), .CI(n29649), .CO(n29651) );
  MXL2HS U32356 ( .A(gray_img[1414]), .B(gray_img[1286]), .S(n29669), .OB(
        n29685) );
  INV1S U32357 ( .I(gray_img[1294]), .O(n29666) );
  INV1S U32358 ( .I(gray_img[1293]), .O(n29664) );
  INV1S U32359 ( .I(gray_img[1291]), .O(n29660) );
  INV1S U32360 ( .I(gray_img[1290]), .O(n29658) );
  FA1S U32361 ( .A(gray_img[1417]), .B(gray_img[1416]), .CI(intadd_65_CI), 
        .CO(n29657) );
  FA1S U32362 ( .A(n29658), .B(gray_img[1418]), .CI(n29657), .CO(n29659) );
  FA1S U32363 ( .A(n29660), .B(gray_img[1419]), .CI(n29659), .CO(n29661) );
  FA1S U32364 ( .A(n29662), .B(gray_img[1420]), .CI(n29661), .CO(n29663) );
  MXL2HS U32365 ( .A(gray_img[1413]), .B(gray_img[1285]), .S(n29669), .OB(
        n29690) );
  MXL2HS U32366 ( .A(gray_img[1412]), .B(gray_img[1284]), .S(n29669), .OB(
        n29695) );
  MXL2HS U32367 ( .A(gray_img[1411]), .B(gray_img[1283]), .S(n29669), .OB(
        n29700) );
  MXL2HS U32368 ( .A(gray_img[1410]), .B(gray_img[1282]), .S(n29669), .OB(
        n29705) );
  MXL2HS U32369 ( .A(gray_img[1408]), .B(gray_img[1280]), .S(n29669), .OB(
        n30000) );
  MXL2HS U32370 ( .A(gray_img[1409]), .B(gray_img[1281]), .S(n29669), .OB(
        n29710) );
  INV1S U32371 ( .I(n29994), .O(n29996) );
  OAI112HS U32372 ( .C1(n29685), .C2(n29999), .A1(n29684), .B1(n29683), .O(
        n13979) );
  OAI112HS U32373 ( .C1(n29690), .C2(n29999), .A1(n29689), .B1(n29688), .O(
        n13980) );
  OAI112HS U32374 ( .C1(n29695), .C2(n29999), .A1(n29694), .B1(n29693), .O(
        n13981) );
  OAI112HS U32375 ( .C1(n29700), .C2(n29999), .A1(n29699), .B1(n29698), .O(
        n13982) );
  OAI112HS U32376 ( .C1(n29705), .C2(n29999), .A1(n29704), .B1(n29703), .O(
        n13983) );
  OAI112HS U32377 ( .C1(n29710), .C2(n29999), .A1(n29709), .B1(n29708), .O(
        n13984) );
  ND2S U32378 ( .I1(n29739), .I2(n29711), .O(n29714) );
  INV1S U32379 ( .I(n29740), .O(n29742) );
  OAI112HS U32380 ( .C1(n29715), .C2(n29745), .A1(n29714), .B1(n29713), .O(
        n14068) );
  ND2S U32381 ( .I1(n29739), .I2(n29716), .O(n29719) );
  MUX2S U32382 ( .A(n15904), .B(n29740), .S(gray_img[516]), .O(n29717) );
  OA12S U32383 ( .B1(n29837), .B2(n29742), .A1(n29717), .O(n29718) );
  OAI112HS U32384 ( .C1(n29720), .C2(n29745), .A1(n29719), .B1(n29718), .O(
        n14069) );
  ND2S U32385 ( .I1(n29739), .I2(n29721), .O(n29724) );
  OAI112HS U32386 ( .C1(n29725), .C2(n29745), .A1(n29724), .B1(n29723), .O(
        n14070) );
  ND2S U32387 ( .I1(n29739), .I2(n29726), .O(n29729) );
  OAI112HS U32388 ( .C1(n29730), .C2(n29745), .A1(n29729), .B1(n29728), .O(
        n14071) );
  MUX2S U32389 ( .A(gray_img[1152]), .B(gray_img[1024]), .S(n29731), .O(n29732) );
  ND2S U32390 ( .I1(n29739), .I2(n29732), .O(n29736) );
  OAI112HS U32391 ( .C1(n29737), .C2(n29745), .A1(n29736), .B1(n29735), .O(
        n13746) );
  ND2S U32392 ( .I1(n29739), .I2(n29738), .O(n29744) );
  OAI112HS U32393 ( .C1(n29746), .C2(n29745), .A1(n29744), .B1(n29743), .O(
        n14072) );
  INV1S U32394 ( .I(gray_img[1298]), .O(n29749) );
  INV1S U32395 ( .I(gray_img[1311]), .O(n29772) );
  INV1S U32396 ( .I(gray_img[1309]), .O(n29768) );
  INV1S U32397 ( .I(gray_img[1307]), .O(n29764) );
  INV1S U32398 ( .I(gray_img[1306]), .O(n29762) );
  INV1S U32399 ( .I(gray_img[1305]), .O(n29760) );
  MXL2HS U32400 ( .A(gray_img[1310]), .B(gray_img[1438]), .S(n29895), .OB(
        n29786) );
  MXL2HS U32401 ( .A(gray_img[1309]), .B(gray_img[1437]), .S(n29895), .OB(
        n29861) );
  MXL2HS U32402 ( .A(gray_img[1308]), .B(gray_img[1436]), .S(n29895), .OB(
        n29866) );
  MXL2HS U32403 ( .A(gray_img[1307]), .B(gray_img[1435]), .S(n29895), .OB(
        n29871) );
  MXL2HS U32404 ( .A(gray_img[1306]), .B(gray_img[1434]), .S(n29895), .OB(
        n29876) );
  MXL2HS U32405 ( .A(gray_img[1305]), .B(gray_img[1433]), .S(n29895), .OB(
        n29891) );
  INV1S U32406 ( .I(n29783), .O(n29782) );
  NR2 U32407 ( .I1(n29680), .I2(n29782), .O(n29904) );
  OR2 U32408 ( .I1(n29680), .I2(n29783), .O(n29894) );
  ND2S U32409 ( .I1(n15890), .I2(n29898), .O(n29784) );
  OAI112HS U32410 ( .C1(n29894), .C2(n29786), .A1(n29785), .B1(n29784), .O(
        n29787) );
  INV1S U32411 ( .I(gray_img[1182]), .O(n29797) );
  INV1S U32412 ( .I(gray_img[1181]), .O(n29795) );
  INV1S U32413 ( .I(gray_img[1180]), .O(n29793) );
  INV1S U32414 ( .I(gray_img[1179]), .O(n29791) );
  MAO222S U32415 ( .A1(gray_img[1048]), .B1(gray_img[1049]), .C1(intadd_86_CI), 
        .O(n29789) );
  FA1S U32416 ( .A(intadd_86_B_1_), .B(gray_img[1050]), .CI(n29789), .CO(
        n29790) );
  FA1S U32417 ( .A(n29791), .B(gray_img[1051]), .CI(n29790), .CO(n29792) );
  FA1S U32418 ( .A(n29793), .B(gray_img[1052]), .CI(n29792), .CO(n29794) );
  MXL2HS U32419 ( .A(gray_img[1182]), .B(gray_img[1054]), .S(n29812), .OB(
        n29828) );
  INV1S U32420 ( .I(gray_img[1174]), .O(n29809) );
  INV1S U32421 ( .I(gray_img[1173]), .O(n29807) );
  INV1S U32422 ( .I(gray_img[1172]), .O(n29805) );
  INV1S U32423 ( .I(gray_img[1169]), .O(n29800) );
  MXL2HS U32424 ( .A(gray_img[1181]), .B(gray_img[1053]), .S(n29812), .OB(
        n29834) );
  MXL2HS U32425 ( .A(gray_img[1180]), .B(gray_img[1052]), .S(n29812), .OB(
        n29840) );
  MXL2HS U32426 ( .A(gray_img[1179]), .B(gray_img[1051]), .S(n29812), .OB(
        n29846) );
  MXL2HS U32427 ( .A(gray_img[1178]), .B(gray_img[1050]), .S(n29812), .OB(
        n29852) );
  MXL2HS U32428 ( .A(gray_img[1176]), .B(gray_img[1048]), .S(n29812), .OB(
        n29858) );
  MXL2HS U32429 ( .A(gray_img[1177]), .B(gray_img[1049]), .S(n29812), .OB(
        n29888) );
  OR2 U32430 ( .I1(n29680), .I2(n29821), .O(n29887) );
  INV1S U32431 ( .I(n29821), .O(n29822) );
  ND2S U32432 ( .I1(n29880), .I2(n29823), .O(n29827) );
  INV1S U32433 ( .I(n29881), .O(n29883) );
  OAI112HS U32434 ( .C1(n29828), .C2(n29887), .A1(n29827), .B1(n29826), .O(
        n14058) );
  ND2S U32435 ( .I1(n29880), .I2(n29829), .O(n29833) );
  OAI112HS U32436 ( .C1(n29834), .C2(n29887), .A1(n29833), .B1(n29832), .O(
        n14059) );
  ND2S U32437 ( .I1(n29880), .I2(n29835), .O(n29839) );
  OAI112HS U32438 ( .C1(n29840), .C2(n29887), .A1(n29839), .B1(n29838), .O(
        n14060) );
  ND2S U32439 ( .I1(n29880), .I2(n29841), .O(n29845) );
  OAI112HS U32440 ( .C1(n29846), .C2(n29887), .A1(n29845), .B1(n29844), .O(
        n14061) );
  ND2S U32441 ( .I1(n29880), .I2(n29847), .O(n29851) );
  OAI112HS U32442 ( .C1(n29852), .C2(n29887), .A1(n29851), .B1(n29850), .O(
        n14062) );
  MUX2S U32443 ( .A(gray_img[1168]), .B(gray_img[1040]), .S(n29853), .O(n29854) );
  ND2S U32444 ( .I1(n29880), .I2(n29854), .O(n29857) );
  OAI112HS U32445 ( .C1(n29858), .C2(n29887), .A1(n29857), .B1(n29856), .O(
        n13745) );
  OAI112HS U32446 ( .C1(n29894), .C2(n29861), .A1(n29860), .B1(n29859), .O(
        n29862) );
  OAI112HS U32447 ( .C1(n29894), .C2(n29866), .A1(n29865), .B1(n29864), .O(
        n29867) );
  OAI112HS U32448 ( .C1(n29894), .C2(n29871), .A1(n29870), .B1(n29869), .O(
        n29872) );
  OAI112HS U32449 ( .C1(n29894), .C2(n29876), .A1(n29875), .B1(n29874), .O(
        n29877) );
  ND2S U32450 ( .I1(n29880), .I2(n29879), .O(n29886) );
  OAI112HS U32451 ( .C1(n29888), .C2(n29887), .A1(n29886), .B1(n29885), .O(
        n14063) );
  OAI112HS U32452 ( .C1(n29894), .C2(n29891), .A1(n29890), .B1(n29889), .O(
        n29892) );
  INV1S U32453 ( .I(n29894), .O(n29897) );
  MUX2S U32454 ( .A(gray_img[1304]), .B(gray_img[1432]), .S(n29895), .O(n29896) );
  ND2S U32455 ( .I1(n29897), .I2(n29896), .O(n29901) );
  ND2S U32456 ( .I1(n15888), .I2(n29898), .O(n29899) );
  ND3S U32457 ( .I1(n29901), .I2(n29900), .I3(n29899), .O(n29902) );
  INV1S U32458 ( .I(gray_img[654]), .O(n29915) );
  INV1S U32459 ( .I(gray_img[653]), .O(n29913) );
  INV1S U32460 ( .I(gray_img[652]), .O(n29911) );
  INV1S U32461 ( .I(gray_img[651]), .O(n29909) );
  INV1S U32462 ( .I(gray_img[650]), .O(n29907) );
  INV1S U32463 ( .I(gray_img[649]), .O(n29905) );
  FA1S U32464 ( .A(gray_img[521]), .B(gray_img[520]), .CI(n29905), .CO(n29906)
         );
  FA1S U32465 ( .A(n29907), .B(gray_img[522]), .CI(n29906), .CO(n29908) );
  FA1S U32466 ( .A(n29909), .B(gray_img[523]), .CI(n29908), .CO(n29910) );
  FA1S U32467 ( .A(n29911), .B(gray_img[524]), .CI(n29910), .CO(n29912) );
  MXL2HS U32468 ( .A(gray_img[518]), .B(gray_img[646]), .S(n30002), .OB(n29943) );
  MXL2HS U32469 ( .A(gray_img[517]), .B(gray_img[645]), .S(n30002), .OB(n29948) );
  MXL2HS U32470 ( .A(gray_img[516]), .B(gray_img[644]), .S(n30002), .OB(n29953) );
  MXL2HS U32471 ( .A(gray_img[515]), .B(gray_img[643]), .S(n30002), .OB(n29958) );
  MXL2HS U32472 ( .A(gray_img[514]), .B(gray_img[642]), .S(n30002), .OB(n29963) );
  MXL2HS U32473 ( .A(gray_img[513]), .B(gray_img[641]), .S(n30002), .OB(n29968) );
  INV1S U32474 ( .I(n29940), .O(n29939) );
  NR2 U32475 ( .I1(n29680), .I2(n29939), .O(n30012) );
  ND2S U32476 ( .I1(n15890), .I2(n30006), .O(n29941) );
  OAI112HS U32477 ( .C1(n30001), .C2(n29943), .A1(n29942), .B1(n29941), .O(
        n29944) );
  OAI112HS U32478 ( .C1(n30001), .C2(n29948), .A1(n29947), .B1(n29946), .O(
        n29949) );
  OAI112HS U32479 ( .C1(n30001), .C2(n29953), .A1(n29952), .B1(n29951), .O(
        n29954) );
  OAI112HS U32480 ( .C1(n30001), .C2(n29958), .A1(n29957), .B1(n29956), .O(
        n29959) );
  OAI112HS U32481 ( .C1(n30001), .C2(n29963), .A1(n29962), .B1(n29961), .O(
        n29964) );
  OAI112HS U32482 ( .C1(n30001), .C2(n29968), .A1(n29967), .B1(n29966), .O(
        n29969) );
  OAI112HS U32483 ( .C1(n30099), .C2(n29973), .A1(n29972), .B1(n29971), .O(
        n29974) );
  OAI112HS U32484 ( .C1(n30099), .C2(n29978), .A1(n29977), .B1(n29976), .O(
        n29979) );
  OAI112HS U32485 ( .C1(n30099), .C2(n29983), .A1(n29982), .B1(n29981), .O(
        n29984) );
  OAI112HS U32486 ( .C1(n30099), .C2(n29988), .A1(n29987), .B1(n29986), .O(
        n29989) );
  MUX2S U32487 ( .A(gray_img[1288]), .B(gray_img[1416]), .S(n29991), .O(n29992) );
  OAI112HS U32488 ( .C1(n30000), .C2(n29999), .A1(n29998), .B1(n29997), .O(
        n13738) );
  INV1S U32489 ( .I(n30001), .O(n30004) );
  MUX2S U32490 ( .A(gray_img[512]), .B(gray_img[640]), .S(n30002), .O(n30003)
         );
  ND2S U32491 ( .I1(n30004), .I2(n30003), .O(n30009) );
  MUX2S U32492 ( .A(n30005), .B(n30006), .S(gray_img[256]), .O(n30008) );
  ND2S U32493 ( .I1(n15888), .I2(n30006), .O(n30007) );
  OAI112HS U32494 ( .C1(n30099), .C2(n30015), .A1(n30014), .B1(n30013), .O(
        n30016) );
  MUX2S U32495 ( .A(gray_img[1960]), .B(gray_img[1832]), .S(n30018), .O(n30019) );
  OAI112HS U32496 ( .C1(n30027), .C2(n30026), .A1(n30025), .B1(n30024), .O(
        n13712) );
  INV1S U32497 ( .I(n30028), .O(n30031) );
  MUX2S U32498 ( .A(gray_img[912]), .B(gray_img[784]), .S(n30029), .O(n30030)
         );
  ND2S U32499 ( .I1(n30031), .I2(n30030), .O(n30035) );
  ND2S U32500 ( .I1(n15888), .I2(n30032), .O(n30033) );
  OAI112HS U32501 ( .C1(n30125), .C2(n30041), .A1(n30040), .B1(n30039), .O(
        n30042) );
  OAI112HS U32502 ( .C1(n30125), .C2(n30047), .A1(n30046), .B1(n30045), .O(
        n30048) );
  OAI112HS U32503 ( .C1(n30125), .C2(n30053), .A1(n30052), .B1(n30051), .O(
        n30054) );
  OAI112HS U32504 ( .C1(n30125), .C2(n30060), .A1(n30059), .B1(n30058), .O(
        n30061) );
  MUX2S U32505 ( .A(n27447), .B(n30063), .S(gray_img[856]), .O(n30064) );
  AO12S U32506 ( .B1(n15888), .B2(n30065), .A1(n30064), .O(n14131) );
  INV1S U32507 ( .I(n30066), .O(n30069) );
  MUX2S U32508 ( .A(gray_img[296]), .B(gray_img[424]), .S(n30067), .O(n30068)
         );
  ND2S U32509 ( .I1(n30069), .I2(n30068), .O(n30073) );
  ND2S U32510 ( .I1(n15888), .I2(n30070), .O(n30071) );
  ND3S U32511 ( .I1(n30073), .I2(n30072), .I3(n30071), .O(n30074) );
  INV1S U32512 ( .I(n30077), .O(n30080) );
  MUX2S U32513 ( .A(gray_img[16]), .B(gray_img[144]), .S(n30078), .O(n30079)
         );
  ND2S U32514 ( .I1(n30080), .I2(n30079), .O(n30084) );
  ND2S U32515 ( .I1(n15888), .I2(n30081), .O(n30082) );
  ND3S U32516 ( .I1(n30084), .I2(n30083), .I3(n30082), .O(n30085) );
  INV1S U32517 ( .I(n30088), .O(n30091) );
  MUX2S U32518 ( .A(gray_img[1792]), .B(gray_img[1920]), .S(n30089), .O(n30090) );
  ND2S U32519 ( .I1(n30091), .I2(n30090), .O(n30095) );
  ND2S U32520 ( .I1(n15888), .I2(n30092), .O(n30093) );
  ND3S U32521 ( .I1(n30095), .I2(n30094), .I3(n30093), .O(n30096) );
  INV1S U32522 ( .I(n30099), .O(n30102) );
  MUX2S U32523 ( .A(gray_img[896]), .B(gray_img[768]), .S(n30100), .O(n30101)
         );
  ND2S U32524 ( .I1(n30102), .I2(n30101), .O(n30106) );
  ND2S U32525 ( .I1(n15888), .I2(n30103), .O(n30104) );
  ND3S U32526 ( .I1(n30106), .I2(n30105), .I3(n30104), .O(n30107) );
  INV1S U32527 ( .I(n30110), .O(n30113) );
  MUX2S U32528 ( .A(gray_img[8]), .B(gray_img[136]), .S(n30111), .O(n30112) );
  ND2S U32529 ( .I1(n30113), .I2(n30112), .O(n30116) );
  OAI112HS U32530 ( .C1(n29734), .C2(n30117), .A1(n30116), .B1(n30115), .O(
        n30118) );
  OAI112HS U32531 ( .C1(n30125), .C2(n30124), .A1(n30123), .B1(n30122), .O(
        n30126) );
  NR2 U32532 ( .I1(cnt_bdyn[2]), .I2(n30302), .O(n30367) );
  NR2 U32533 ( .I1(n30387), .I2(n30390), .O(n30393) );
  NR3 U32534 ( .I1(cnt_bdyn[3]), .I2(cnt_bdyn[8]), .I3(n30129), .O(n30130) );
  NR2 U32535 ( .I1(n30222), .I2(n30131), .O(n30134) );
  NR2 U32536 ( .I1(n30452), .I2(n30131), .O(n30133) );
  INV1S U32537 ( .I(n30299), .O(n30221) );
  NR2 U32538 ( .I1(n30221), .I2(n30131), .O(n30136) );
  INV1S U32539 ( .I(cro_mac[13]), .O(n30151) );
  XNR2HS U32540 ( .I1(n30149), .I2(n30148), .O(n30150) );
  MOAI1S U32541 ( .A1(n30220), .A2(n30151), .B1(n30150), .B2(n30218), .O(
        n13598) );
  INV1S U32542 ( .I(cro_mac[10]), .O(n30160) );
  INV1S U32543 ( .I(n30152), .O(n30154) );
  ND2S U32544 ( .I1(n30154), .I2(n30153), .O(n30158) );
  INV1S U32545 ( .I(n30155), .O(n30162) );
  INV1S U32546 ( .I(n30161), .O(n30156) );
  AOI12HS U32547 ( .B1(n30163), .B2(n30162), .A1(n30156), .O(n30157) );
  XOR2HS U32548 ( .I1(n30158), .I2(n30157), .O(n30159) );
  MOAI1S U32549 ( .A1(n30220), .A2(n30160), .B1(n30159), .B2(n30218), .O(
        n13601) );
  INV1S U32550 ( .I(cro_mac[9]), .O(n30166) );
  XNR2HS U32551 ( .I1(n30164), .I2(n30163), .O(n30165) );
  MOAI1S U32552 ( .A1(n30220), .A2(n30166), .B1(n30165), .B2(n30218), .O(
        n13602) );
  INV1S U32553 ( .I(cro_mac[8]), .O(n30174) );
  INV1S U32554 ( .I(n30167), .O(n30169) );
  INV1S U32555 ( .I(n30170), .O(n30179) );
  OAI12HS U32556 ( .B1(n30175), .B2(n30179), .A1(n30176), .O(n30171) );
  XNR2HS U32557 ( .I1(n30172), .I2(n30171), .O(n30173) );
  MOAI1S U32558 ( .A1(n30220), .A2(n30174), .B1(n30173), .B2(n30218), .O(
        n13603) );
  INV1S U32559 ( .I(cro_mac[7]), .O(n30181) );
  INV1S U32560 ( .I(n30175), .O(n30177) );
  XOR2HS U32561 ( .I1(n30179), .I2(n30178), .O(n30180) );
  MOAI1S U32562 ( .A1(n30220), .A2(n30181), .B1(n30180), .B2(n30218), .O(
        n13604) );
  INV1S U32563 ( .I(cro_mac[6]), .O(n30279) );
  INV1S U32564 ( .I(n30182), .O(n30184) );
  XOR2HS U32565 ( .I1(n30186), .I2(n30185), .O(n30187) );
  MOAI1S U32566 ( .A1(n30220), .A2(n30279), .B1(n30187), .B2(n30218), .O(
        n13605) );
  INV1S U32567 ( .I(cro_mac[5]), .O(n30278) );
  XNR2HS U32568 ( .I1(n30191), .I2(n30190), .O(n30192) );
  MOAI1S U32569 ( .A1(n30220), .A2(n30278), .B1(n30192), .B2(n30218), .O(
        n13606) );
  INV1S U32570 ( .I(cro_mac[4]), .O(n30277) );
  INV1S U32571 ( .I(n30193), .O(n30195) );
  XOR2HS U32572 ( .I1(n30197), .I2(n30196), .O(n30198) );
  MOAI1S U32573 ( .A1(n30220), .A2(n30277), .B1(n30198), .B2(n30218), .O(
        n13607) );
  INV1S U32574 ( .I(cro_mac[3]), .O(n30276) );
  INV1S U32575 ( .I(n30199), .O(n30201) );
  ND2S U32576 ( .I1(n30201), .I2(n30200), .O(n30202) );
  XOR2HS U32577 ( .I1(n30203), .I2(n30202), .O(n30204) );
  MOAI1S U32578 ( .A1(n30220), .A2(n30276), .B1(n30204), .B2(n30218), .O(
        n13608) );
  INV1S U32579 ( .I(cro_mac[2]), .O(n30275) );
  ND2S U32580 ( .I1(n30206), .I2(n30205), .O(n30207) );
  XNR2HS U32581 ( .I1(n30208), .I2(n30207), .O(n30209) );
  MOAI1S U32582 ( .A1(n30220), .A2(n30275), .B1(n30209), .B2(n30218), .O(
        n13609) );
  INV1S U32583 ( .I(cro_mac[1]), .O(n30274) );
  INV1S U32584 ( .I(n30210), .O(n30212) );
  ND2S U32585 ( .I1(n30212), .I2(n30211), .O(n30213) );
  XOR2HS U32586 ( .I1(n30216), .I2(n30213), .O(n30214) );
  MOAI1S U32587 ( .A1(n30220), .A2(n30274), .B1(n30214), .B2(n30218), .O(
        n13610) );
  INV1S U32588 ( .I(cro_mac[0]), .O(n30273) );
  OR2S U32589 ( .I1(cro_mac[0]), .I2(n30215), .O(n30217) );
  AN2S U32590 ( .I1(n30217), .I2(n30216), .O(n30219) );
  MOAI1S U32591 ( .A1(n30220), .A2(n30273), .B1(n30219), .B2(n30218), .O(
        n13611) );
  MOAI1S U32592 ( .A1(n30338), .A2(n30452), .B1(C551_DATA2_4), .B2(n30349), 
        .O(gray_scale_2_n[4]) );
  MOAI1S U32593 ( .A1(n30421), .A2(n30452), .B1(C551_DATA2_3), .B2(n30349), 
        .O(gray_scale_2_n[3]) );
  MOAI1S U32594 ( .A1(n30418), .A2(n30452), .B1(C551_DATA2_2), .B2(n30349), 
        .O(gray_scale_2_n[2]) );
  MOAI1S U32595 ( .A1(n30417), .A2(n30452), .B1(C551_DATA2_1), .B2(n30349), 
        .O(gray_scale_2_n[1]) );
  MOAI1S U32596 ( .A1(n30416), .A2(n30452), .B1(C551_DATA2_0), .B2(n30349), 
        .O(gray_scale_2_n[0]) );
  NR2 U32597 ( .I1(n30221), .I2(n30423), .O(C1_Z_6) );
  MOAI1S U32598 ( .A1(n30423), .A2(n30222), .B1(image[6]), .B2(n30299), .O(
        C1_Z_5) );
  MOAI1S U32599 ( .A1(n30338), .A2(n30222), .B1(image[5]), .B2(n30299), .O(
        C1_Z_4) );
  MOAI1S U32600 ( .A1(n30421), .A2(n30222), .B1(image[4]), .B2(n30299), .O(
        C1_Z_3) );
  MOAI1S U32601 ( .A1(n30418), .A2(n30222), .B1(image[3]), .B2(n30299), .O(
        C1_Z_2) );
  MOAI1S U32602 ( .A1(n30417), .A2(n30222), .B1(image[2]), .B2(n30299), .O(
        C1_Z_1) );
  MOAI1S U32603 ( .A1(n30416), .A2(n30222), .B1(image[1]), .B2(n30299), .O(
        C1_Z_0) );
  XOR2HS U32604 ( .I1(gray_scale_2[7]), .I2(DP_OP_989J1_126_3015_n1), .O(
        n30223) );
  NR2 U32605 ( .I1(cnt_20[5]), .I2(cnt_20[4]), .O(n30225) );
  NR2 U32606 ( .I1(cnt_20[1]), .I2(cnt_20[2]), .O(n30224) );
  AN4S U32607 ( .I1(n30225), .I2(cnt_20[3]), .I3(n30224), .I4(cnt_20[0]), .O(
        n30380) );
  MUX2S U32608 ( .A(cro_mac[7]), .B(cro_mac_store[6]), .S(n30226), .O(N7773)
         );
  MUX2S U32609 ( .A(cro_mac[8]), .B(cro_mac_store[7]), .S(n30226), .O(N7774)
         );
  MUX2S U32610 ( .A(cro_mac[9]), .B(cro_mac_store[8]), .S(n30226), .O(N7775)
         );
  MUX2S U32611 ( .A(cro_mac[10]), .B(cro_mac_store[9]), .S(n30226), .O(N7776)
         );
  MUX2S U32612 ( .A(cro_mac[11]), .B(cro_mac_store[10]), .S(n30226), .O(N7777)
         );
  MUX2S U32613 ( .A(cro_mac[12]), .B(cro_mac_store[11]), .S(n30226), .O(N7778)
         );
  MUX2S U32614 ( .A(cro_mac[13]), .B(cro_mac_store[12]), .S(n30226), .O(N7779)
         );
  MUX2S U32615 ( .A(cro_mac[14]), .B(cro_mac_store[13]), .S(n30226), .O(N7780)
         );
  MUX2S U32616 ( .A(cro_mac[15]), .B(cro_mac_store[14]), .S(n30226), .O(N7781)
         );
  MUX2S U32617 ( .A(cro_mac[16]), .B(cro_mac_store[15]), .S(n30226), .O(N7782)
         );
  MUX2S U32618 ( .A(cro_mac[17]), .B(cro_mac_store[16]), .S(n30226), .O(N7783)
         );
  MUX2S U32619 ( .A(cro_mac[18]), .B(cro_mac_store[17]), .S(n30226), .O(N7784)
         );
  MUX2S U32620 ( .A(cro_mac[19]), .B(cro_mac_store[18]), .S(n30226), .O(N7785)
         );
  AN2S U32621 ( .I1(out_valid_a1), .I2(cro_mac_store[19]), .O(out_value_a1) );
  NR2 U32622 ( .I1(cnt_20[0]), .I2(n30360), .O(cnt_20_n[0]) );
  INV1S U32623 ( .I(n30227), .O(n30229) );
  AN2S U32624 ( .I1(cnt_20[2]), .I2(n30229), .O(n30231) );
  NR3 U32625 ( .I1(cnt_20[5]), .I2(cnt_20[3]), .I3(cnt_20[2]), .O(n30228) );
  AO13S U32626 ( .B1(n30229), .B2(cnt_20[4]), .B3(n30228), .A1(n30360), .O(
        n30237) );
  NR2 U32627 ( .I1(cnt_20[2]), .I2(n30229), .O(n30230) );
  NR3 U32628 ( .I1(n30231), .I2(n30237), .I3(n30230), .O(cnt_20_n[2]) );
  AN2S U32629 ( .I1(cnt_20[3]), .I2(n30231), .O(n30233) );
  NR2 U32630 ( .I1(cnt_20[3]), .I2(n30231), .O(n30232) );
  NR3 U32631 ( .I1(n30233), .I2(n30237), .I3(n30232), .O(cnt_20_n[3]) );
  AN2S U32632 ( .I1(cnt_20[4]), .I2(n30233), .O(n30235) );
  NR2 U32633 ( .I1(cnt_20[4]), .I2(n30233), .O(n30234) );
  NR3 U32634 ( .I1(n30235), .I2(n30237), .I3(n30234), .O(cnt_20_n[4]) );
  MOAI1S U32635 ( .A1(cnt_20[5]), .A2(n30235), .B1(cnt_20[5]), .B2(n30235), 
        .O(n30236) );
  NR2 U32636 ( .I1(n30237), .I2(n30236), .O(cnt_20_n[5]) );
  INV1S U32637 ( .I(n30238), .O(n30240) );
  ND2S U32638 ( .I1(n30240), .I2(n30239), .O(n30426) );
  AO12S U32639 ( .B1(n30242), .B2(n30241), .A1(n30426), .O(n30249) );
  NR2 U32640 ( .I1(medfilt_cnt[0]), .I2(n30249), .O(N7502) );
  MOAI1S U32641 ( .A1(medfilt_cnt[1]), .A2(medfilt_cnt[0]), .B1(medfilt_cnt[1]), .B2(medfilt_cnt[0]), .O(n30243) );
  NR2 U32642 ( .I1(n30249), .I2(n30243), .O(N7503) );
  ND2S U32643 ( .I1(medfilt_cnt[1]), .I2(medfilt_cnt[0]), .O(n30245) );
  MOAI1S U32644 ( .A1(n30246), .A2(n30245), .B1(n30246), .B2(n30245), .O(
        n30244) );
  NR2 U32645 ( .I1(n30249), .I2(n30244), .O(N7504) );
  NR2 U32646 ( .I1(n30246), .I2(n30245), .O(n30247) );
  MOAI1S U32647 ( .A1(medfilt_cnt[3]), .A2(n30247), .B1(medfilt_cnt[3]), .B2(
        n30247), .O(n30248) );
  NR2 U32648 ( .I1(n30249), .I2(n30248), .O(N7505) );
  MOAI1S U32649 ( .A1(n30305), .A2(n30251), .B1(n30305), .B2(n30251), .O(
        n30250) );
  NR2 U32650 ( .I1(n30254), .I2(n30250), .O(cnt_dyn_n[2]) );
  NR2 U32651 ( .I1(n30305), .I2(n30251), .O(n30252) );
  MOAI1S U32652 ( .A1(cnt_dyn[3]), .A2(n30252), .B1(cnt_dyn[3]), .B2(n30252), 
        .O(n30253) );
  NR2 U32653 ( .I1(n30254), .I2(n30253), .O(cnt_dyn_n[3]) );
  INV1S U32654 ( .I(n30255), .O(n30256) );
  OAI12HS U32655 ( .B1(last_in_valid2), .B2(n30257), .A1(n30256), .O(n30272)
         );
  NR2 U32656 ( .I1(cnt[0]), .I2(n30272), .O(cnt_n[0]) );
  ND2S U32657 ( .I1(cnt[0]), .I2(cnt[1]), .O(n30258) );
  INV1S U32658 ( .I(n30258), .O(n30260) );
  NR2 U32659 ( .I1(cnt[0]), .I2(cnt[1]), .O(n30428) );
  NR3 U32660 ( .I1(n30260), .I2(n30428), .I3(n30272), .O(cnt_n[1]) );
  NR2 U32661 ( .I1(n30259), .I2(n30258), .O(n30262) );
  NR2 U32662 ( .I1(cnt[2]), .I2(n30260), .O(n30261) );
  NR3 U32663 ( .I1(n30262), .I2(n30272), .I3(n30261), .O(cnt_n[2]) );
  AN2S U32664 ( .I1(cnt[3]), .I2(n30262), .O(n30264) );
  NR2 U32665 ( .I1(cnt[3]), .I2(n30262), .O(n30263) );
  NR3 U32666 ( .I1(n30264), .I2(n30272), .I3(n30263), .O(cnt_n[3]) );
  AN2S U32667 ( .I1(cnt[4]), .I2(n30264), .O(n30266) );
  NR2 U32668 ( .I1(cnt[4]), .I2(n30264), .O(n30265) );
  NR3 U32669 ( .I1(n30266), .I2(n30272), .I3(n30265), .O(cnt_n[4]) );
  AN2S U32670 ( .I1(cnt[5]), .I2(n30266), .O(n30268) );
  NR2 U32671 ( .I1(cnt[5]), .I2(n30266), .O(n30267) );
  NR3 U32672 ( .I1(n30268), .I2(n30272), .I3(n30267), .O(cnt_n[5]) );
  AN2S U32673 ( .I1(cnt[6]), .I2(n30268), .O(n30270) );
  NR2 U32674 ( .I1(cnt[6]), .I2(n30268), .O(n30269) );
  NR3 U32675 ( .I1(n30270), .I2(n30272), .I3(n30269), .O(cnt_n[6]) );
  MOAI1S U32676 ( .A1(cnt[7]), .A2(n30270), .B1(cnt[7]), .B2(n30270), .O(
        n30271) );
  NR2 U32677 ( .I1(n30272), .I2(n30271), .O(cnt_n[7]) );
  NR2 U32678 ( .I1(n30226), .I2(n30273), .O(N7766) );
  MOAI1S U32679 ( .A1(n30226), .A2(n30274), .B1(n30226), .B2(cro_mac_store[0]), 
        .O(N7767) );
  MOAI1S U32680 ( .A1(n30226), .A2(n30275), .B1(n30226), .B2(cro_mac_store[1]), 
        .O(N7768) );
  MOAI1S U32681 ( .A1(n30226), .A2(n30276), .B1(n30226), .B2(cro_mac_store[2]), 
        .O(N7769) );
  MOAI1S U32682 ( .A1(n30226), .A2(n30277), .B1(n30226), .B2(cro_mac_store[3]), 
        .O(N7770) );
  MOAI1S U32683 ( .A1(n30226), .A2(n30278), .B1(n30226), .B2(cro_mac_store[4]), 
        .O(N7771) );
  MOAI1S U32684 ( .A1(n30226), .A2(n30279), .B1(n30226), .B2(cro_mac_store[5]), 
        .O(N7772) );
  INV1S U32685 ( .I(image_size_reg_master[0]), .O(n30395) );
  ND2S U32686 ( .I1(image_size_reg_master[1]), .I2(n30395), .O(n30319) );
  ND2S U32687 ( .I1(image_size_reg_master[0]), .I2(n30394), .O(n30318) );
  INV1S U32688 ( .I(cnt_bdyn[4]), .O(n30313) );
  NR2 U32689 ( .I1(image_size_reg_master[0]), .I2(image_size_reg_master[1]), 
        .O(n30311) );
  INV1S U32690 ( .I(n30311), .O(n30316) );
  OA222S U32691 ( .A1(n30280), .A2(n30319), .B1(n30323), .B2(n30318), .C1(
        n30313), .C2(n30316), .O(n30282) );
  NR2 U32692 ( .I1(n30282), .I2(n30281), .O(n30283) );
  ND2S U32693 ( .I1(image_size_reg_master[0]), .I2(image_size_reg_master[1]), 
        .O(n30301) );
  AOI22S U32694 ( .A1(n30451), .A2(n30283), .B1(mem_we_a_reg), .B2(n30301), 
        .O(n30284) );
  NR2 U32695 ( .I1(n30284), .I2(n30390), .O(N442) );
  OR2B1S U32696 ( .I1(cs_d1[1]), .B1(n30290), .O(n30334) );
  INV1S U32697 ( .I(n30334), .O(n30329) );
  AO222S U32698 ( .A1(n30451), .A2(gray_scale_2_s[0]), .B1(n30298), .B2(
        gray_scale_1_s[0]), .C1(n30299), .C2(gray_scale_0_s[0]), .O(n30291) );
  AN2S U32699 ( .I1(n30329), .I2(n30291), .O(mem_data_a_in[0]) );
  AO222S U32700 ( .A1(n30451), .A2(gray_scale_2_s[1]), .B1(n30298), .B2(
        gray_scale_1_s[1]), .C1(n30299), .C2(gray_scale_0_s[1]), .O(n30292) );
  AN2S U32701 ( .I1(n30329), .I2(n30292), .O(mem_data_a_in[1]) );
  AO222S U32702 ( .A1(n30451), .A2(gray_scale_2_s[2]), .B1(n30298), .B2(
        gray_scale_1_s[2]), .C1(n30299), .C2(gray_scale_0_s[2]), .O(n30293) );
  AN2S U32703 ( .I1(n30329), .I2(n30293), .O(mem_data_a_in[2]) );
  AO222S U32704 ( .A1(n30451), .A2(gray_scale_2_s[3]), .B1(n30298), .B2(
        gray_scale_1_s[3]), .C1(n30299), .C2(gray_scale_0_s[3]), .O(n30294) );
  AN2S U32705 ( .I1(n30329), .I2(n30294), .O(mem_data_a_in[3]) );
  AO222S U32706 ( .A1(n30451), .A2(gray_scale_2_s[4]), .B1(n30298), .B2(
        gray_scale_1_s[4]), .C1(n30299), .C2(gray_scale_0_s[4]), .O(n30295) );
  AN2S U32707 ( .I1(n30329), .I2(n30295), .O(mem_data_a_in[4]) );
  AO222S U32708 ( .A1(n30451), .A2(gray_scale_2_s[5]), .B1(n30299), .B2(
        gray_scale_0_s[5]), .C1(n30298), .C2(gray_scale_1_s[5]), .O(n30296) );
  AN2S U32709 ( .I1(n30329), .I2(n30296), .O(mem_data_a_in[5]) );
  AO222S U32710 ( .A1(n30451), .A2(gray_scale_2_s[6]), .B1(n30299), .B2(
        gray_scale_0_s[6]), .C1(n30298), .C2(gray_scale_1_s[6]), .O(n30297) );
  AN2S U32711 ( .I1(n30329), .I2(n30297), .O(mem_data_a_in[6]) );
  AO222S U32712 ( .A1(n30451), .A2(gray_scale_2_s[7]), .B1(n30299), .B2(
        gray_scale_0_s[7]), .C1(gray_scale_1_s[7]), .C2(n30298), .O(n30300) );
  AN2S U32713 ( .I1(n30329), .I2(n30300), .O(mem_data_a_in[7]) );
  OR2S U32714 ( .I1(mem_we_a_reg), .I2(n30334), .O(mem_we_a) );
  OAI22S U32715 ( .A1(cnt_bdyn[0]), .A2(n30335), .B1(n30333), .B2(n30329), .O(
        mem_addr_a[0]) );
  NR2 U32716 ( .I1(n30302), .I2(n30303), .O(n30368) );
  OAI22S U32717 ( .A1(n30368), .A2(n30335), .B1(n30349), .B2(n30329), .O(
        mem_addr_a[1]) );
  NR2 U32718 ( .I1(n30311), .I2(n30335), .O(n30304) );
  MOAI1S U32719 ( .A1(n30303), .A2(n30365), .B1(n30303), .B2(n30365), .O(
        n30310) );
  MOAI1S U32720 ( .A1(n30329), .A2(n30305), .B1(n30304), .B2(n30310), .O(
        mem_addr_a[2]) );
  MOAI1S U32721 ( .A1(n30330), .A2(n30306), .B1(n30330), .B2(n30306), .O(
        n30315) );
  OR2S U32722 ( .I1(n30334), .I2(n30319), .O(n30332) );
  OAI22S U32723 ( .A1(n30315), .A2(n30332), .B1(n30307), .B2(n30329), .O(
        mem_addr_a[3]) );
  MOAI1S U32724 ( .A1(n30308), .A2(n30313), .B1(n30308), .B2(n30313), .O(
        n30317) );
  OR2S U32725 ( .I1(n30334), .I2(n30318), .O(n30325) );
  OAI22S U32726 ( .A1(n30315), .A2(n30325), .B1(n30372), .B2(n30329), .O(
        n30309) );
  AOI13HS U32727 ( .B1(n30329), .B2(n30311), .B3(n30310), .A1(n30309), .O(
        n30312) );
  OAI12HS U32728 ( .B1(n30317), .B2(n30332), .A1(n30312), .O(mem_addr_a[4]) );
  ND2S U32729 ( .I1(n30322), .I2(n30313), .O(n30314) );
  AOI22S U32730 ( .A1(n30322), .A2(n30321), .B1(cnt_bdyn[5]), .B2(n30314), .O(
        n30324) );
  OA222S U32731 ( .A1(n30319), .A2(n30324), .B1(n30318), .B2(n30317), .C1(
        n30316), .C2(n30315), .O(n30320) );
  OAI22S U32732 ( .A1(n30334), .A2(n30320), .B1(n30329), .B2(n30369), .O(
        mem_addr_a[5]) );
  ND2S U32733 ( .I1(n30322), .I2(n30321), .O(n30327) );
  MOAI1S U32734 ( .A1(n30323), .A2(n30327), .B1(n30323), .B2(n30327), .O(
        n30326) );
  OAI222S U32735 ( .A1(n30332), .A2(n30326), .B1(n30325), .B2(n30324), .C1(
        n30365), .C2(n30329), .O(mem_addr_a[6]) );
  NR2 U32736 ( .I1(cnt_bdyn[6]), .I2(n30327), .O(n30328) );
  MOAI1S U32737 ( .A1(cnt_bdyn[7]), .A2(n30328), .B1(cnt_bdyn[7]), .B2(n30328), 
        .O(n30331) );
  OAI22S U32738 ( .A1(n30332), .A2(n30331), .B1(n30330), .B2(n30329), .O(
        mem_addr_a[7]) );
  MOAI1S U32739 ( .A1(n30333), .A2(n30335), .B1(read_layer[0]), .B2(n30334), 
        .O(mem_addr_a[8]) );
  MOAI1S U32740 ( .A1(n30349), .A2(n30335), .B1(read_layer[1]), .B2(n30334), 
        .O(mem_addr_a[9]) );
  MOAI1S U32741 ( .A1(n30338), .A2(n30452), .B1(n30337), .B2(n30349), .O(
        n15822) );
  MOAI1S U32742 ( .A1(n30421), .A2(n30452), .B1(n30340), .B2(n30349), .O(
        n15821) );
  MOAI1S U32743 ( .A1(n30418), .A2(n30452), .B1(n30342), .B2(n30349), .O(
        n15820) );
  MOAI1S U32744 ( .A1(n30417), .A2(n30452), .B1(n30344), .B2(n30349), .O(
        n15819) );
  MOAI1S U32745 ( .A1(n30416), .A2(n30452), .B1(n30346), .B2(n30349), .O(
        n15818) );
  MOAI1S U32746 ( .A1(n30415), .A2(n30452), .B1(n30348), .B2(n30349), .O(
        n15817) );
  INV1S U32747 ( .I(image[0]), .O(n30414) );
  MOAI1S U32748 ( .A1(n30414), .A2(n30452), .B1(n30350), .B2(n30349), .O(
        n15816) );
  NR2 U32749 ( .I1(n30353), .I2(n30352), .O(n30355) );
  MOAI1S U32750 ( .A1(cnt_bdyn[8]), .A2(n30355), .B1(cnt_bdyn[8]), .B2(n30355), 
        .O(n30351) );
  NR2 U32751 ( .I1(n30360), .I2(n30351), .O(n15804) );
  AN2S U32752 ( .I1(n30353), .I2(n30352), .O(n30354) );
  NR3 U32753 ( .I1(n30355), .I2(n30360), .I3(n30354), .O(n15803) );
  NR2 U32754 ( .I1(cnt_bdyn[5]), .I2(n30356), .O(n30357) );
  NR3 U32755 ( .I1(n30358), .I2(n30360), .I3(n30357), .O(n15801) );
  NR2 U32756 ( .I1(n30360), .I2(n30359), .O(n30370) );
  ND2S U32757 ( .I1(n30371), .I2(n30363), .O(n30362) );
  MOAI1S U32758 ( .A1(n30364), .A2(n30363), .B1(cnt_bdyn[3]), .B2(n30362), .O(
        n15799) );
  ND2S U32759 ( .I1(n30370), .I2(n30364), .O(n30366) );
  OAI22S U32760 ( .A1(n30367), .A2(n30366), .B1(n30365), .B2(n30371), .O(
        n15798) );
  MOAI1S U32761 ( .A1(n30369), .A2(n30371), .B1(n30370), .B2(n30368), .O(
        n15797) );
  MOAI1S U32762 ( .A1(n30372), .A2(n30371), .B1(n30372), .B2(n30370), .O(
        n15796) );
  NR2 U32763 ( .I1(action_done), .I2(n30432), .O(n30385) );
  AN4B1S U32764 ( .I1(n30374), .I2(n30373), .I3(cnt_cro_x[0]), .B1(
        cnt_cro_y[3]), .O(n30377) );
  NR2 U32765 ( .I1(cnt_cro_y[1]), .I2(cnt_cro_x[2]), .O(n30376) );
  AN4B1S U32766 ( .I1(n30377), .I2(n30376), .I3(n30375), .B1(cnt_cro_y[2]), 
        .O(n30378) );
  ND3S U32767 ( .I1(n30380), .I2(n30379), .I3(n30378), .O(n30434) );
  AN4B1S U32768 ( .I1(out_valid), .I2(set_cnt[1]), .I3(set_cnt[2]), .B1(n30434), .O(n30381) );
  ND2S U32769 ( .I1(set_cnt[0]), .I2(n30381), .O(n30382) );
  AO13S U32770 ( .B1(n30383), .B2(n30385), .B3(n30382), .A1(n30411), .O(n15794) );
  NR2 U32771 ( .I1(n30385), .I2(n30384), .O(n30386) );
  AOI13HS U32772 ( .B1(n30388), .B2(in_valid2), .B3(n30387), .A1(n30386), .O(
        n30392) );
  AOI13HS U32773 ( .B1(n30392), .B2(n30391), .B3(n30390), .A1(n30389), .O(
        n15792) );
  AN2B1S U32774 ( .I1(n30393), .B1(last_in_valid_d1), .O(n30396) );
  MOAI1S U32775 ( .A1(n30396), .A2(n30394), .B1(n30396), .B2(
        image_size_in_reg[1]), .O(n15791) );
  MOAI1S U32776 ( .A1(n30396), .A2(n30395), .B1(n30396), .B2(
        image_size_in_reg[0]), .O(n15790) );
  AO12S U32777 ( .B1(cnt[1]), .B2(cnt[2]), .A1(n30397), .O(n30399) );
  OR2B1S U32778 ( .I1(n30398), .B1(n30399), .O(n30405) );
  MOAI1S U32779 ( .A1(n30405), .A2(n30401), .B1(n30405), .B2(action_reg[21]), 
        .O(n15788) );
  OR2B1S U32780 ( .I1(n30400), .B1(n30399), .O(n30407) );
  MOAI1S U32781 ( .A1(n30407), .A2(n30401), .B1(n30407), .B2(action_reg[18]), 
        .O(n30402) );
  AO12S U32782 ( .B1(n18401), .B2(action_reg[21]), .A1(n30402), .O(n15787) );
  MOAI1S U32783 ( .A1(n30405), .A2(n30403), .B1(n30405), .B2(action_reg[22]), 
        .O(n15780) );
  MOAI1S U32784 ( .A1(n30407), .A2(n30403), .B1(n30407), .B2(action_reg[19]), 
        .O(n30404) );
  AO12S U32785 ( .B1(n18401), .B2(action_reg[22]), .A1(n30404), .O(n15779) );
  MOAI1S U32786 ( .A1(n30405), .A2(n30406), .B1(n30405), .B2(action_reg[23]), 
        .O(n15772) );
  MOAI1S U32787 ( .A1(n30407), .A2(n30406), .B1(n30407), .B2(action_reg[20]), 
        .O(n30408) );
  AO12S U32788 ( .B1(n18401), .B2(action_reg[23]), .A1(n30408), .O(n15771) );
  MOAI1S U32789 ( .A1(n30409), .A2(n30412), .B1(n30411), .B2(action_reg[0]), 
        .O(n15760) );
  MOAI1S U32790 ( .A1(n30410), .A2(n30412), .B1(n30411), .B2(action_reg[1]), 
        .O(n15759) );
  MOAI1S U32791 ( .A1(n30413), .A2(n30412), .B1(n30411), .B2(action_reg[2]), 
        .O(n15758) );
  MOAI1S U32792 ( .A1(n30414), .A2(n30420), .B1(gray_scale_0[0]), .B2(n30419), 
        .O(n15744) );
  MOAI1S U32793 ( .A1(n30415), .A2(n30420), .B1(gray_scale_0[1]), .B2(n30419), 
        .O(n15743) );
  MOAI1S U32794 ( .A1(n30416), .A2(n30420), .B1(gray_scale_0[2]), .B2(n30419), 
        .O(n15742) );
  MOAI1S U32795 ( .A1(n30417), .A2(n30420), .B1(gray_scale_0[3]), .B2(n30419), 
        .O(n15741) );
  MOAI1S U32796 ( .A1(n30418), .A2(n30420), .B1(gray_scale_0[4]), .B2(n30419), 
        .O(n15740) );
  MOAI1S U32797 ( .A1(n30421), .A2(n30420), .B1(gray_scale_0[5]), .B2(n30419), 
        .O(n15739) );
  MOAI1S U32798 ( .A1(n30424), .A2(n30423), .B1(n30422), .B2(gray_scale_0[7]), 
        .O(n15737) );
  MOAI1S U32799 ( .A1(n30427), .A2(n30426), .B1(n30427), .B2(n30425), .O(
        n15736) );
  AN4B1S U32800 ( .I1(n30429), .I2(last_in_valid2), .I3(n30428), .B1(cnt[2]), 
        .O(n30430) );
  MUX2S U32801 ( .A(read_layer[1]), .B(action_in_reg[1]), .S(n30430), .O(
        n13590) );
  MUX2S U32802 ( .A(read_layer[0]), .B(action_in_reg[0]), .S(n30430), .O(
        n13589) );
  ND2S U32803 ( .I1(n30432), .I2(set_cnt[0]), .O(n30431) );
  OA12S U32804 ( .B1(n30432), .B2(set_cnt[0]), .A1(n30431), .O(n13588) );
  MOAI1S U32805 ( .A1(set_cnt[1]), .A2(n30431), .B1(set_cnt[1]), .B2(n30431), 
        .O(n13587) );
  ND3S U32806 ( .I1(n30432), .I2(set_cnt[0]), .I3(set_cnt[1]), .O(n30433) );
  MOAI1S U32807 ( .A1(set_cnt[2]), .A2(n30433), .B1(set_cnt[2]), .B2(n30433), 
        .O(n13586) );
  MOAI1S U32808 ( .A1(out_valid_a1), .A2(n30434), .B1(out_valid_a1), .B2(
        n30434), .O(n13585) );
  MUX2S U32809 ( .A(gray_scale_2[7]), .B(gray_scale_2_s[7]), .S(n30452), .O(
        n13584) );
  AO112S U32810 ( .C1(n30436), .C2(gray_scale_1[1]), .A1(n30435), .B1(n30452), 
        .O(n30437) );
  OA12S U32811 ( .B1(n30451), .B2(gray_scale_1_s[1]), .A1(n30437), .O(n13582)
         );
  OA12S U32812 ( .B1(n30440), .B2(n30439), .A1(n30438), .O(n30441) );
  MOAI1S U32813 ( .A1(n30452), .A2(n30441), .B1(n30452), .B2(gray_scale_1_s[2]), .O(n13581) );
  MUX2S U32814 ( .A(n30442), .B(gray_scale_1_s[3]), .S(n30452), .O(n13580) );
  MOAI1S U32815 ( .A1(n30452), .A2(n30443), .B1(n30452), .B2(gray_scale_1_s[4]), .O(n13579) );
  MUX2S U32816 ( .A(n30444), .B(gray_scale_1_s[5]), .S(n30452), .O(n13578) );
  OA12S U32817 ( .B1(n30447), .B2(n30446), .A1(n30445), .O(n30448) );
  MOAI1S U32818 ( .A1(n30452), .A2(n30448), .B1(n30452), .B2(gray_scale_1_s[6]), .O(n13577) );
  OA222S U32819 ( .A1(n30452), .A2(n30450), .B1(n30452), .B2(n30449), .C1(
        gray_scale_1_s[7]), .C2(n30451), .O(n13576) );
  AO22S U32820 ( .A1(n30452), .A2(gray_scale_0_s[0]), .B1(n30451), .B2(
        gray_scale_0[0]), .O(n13575) );
  AO22S U32821 ( .A1(n30452), .A2(gray_scale_0_s[1]), .B1(n30451), .B2(
        gray_scale_0[1]), .O(n13574) );
  AO22S U32822 ( .A1(n30452), .A2(gray_scale_0_s[2]), .B1(n30451), .B2(
        gray_scale_0[2]), .O(n13573) );
  AO22S U32823 ( .A1(n30452), .A2(gray_scale_0_s[3]), .B1(n30451), .B2(
        gray_scale_0[3]), .O(n13572) );
  AO22S U32824 ( .A1(n30452), .A2(gray_scale_0_s[4]), .B1(n30451), .B2(
        gray_scale_0[4]), .O(n13571) );
  AO22S U32825 ( .A1(n30452), .A2(gray_scale_0_s[5]), .B1(n30451), .B2(
        gray_scale_0[5]), .O(n13570) );
  AO22S U32826 ( .A1(n30452), .A2(gray_scale_0_s[6]), .B1(n30451), .B2(
        gray_scale_0[6]), .O(n13569) );
  AO22S U32827 ( .A1(n30452), .A2(gray_scale_0_s[7]), .B1(n30451), .B2(
        gray_scale_0[7]), .O(n13568) );
  MUX2S U32828 ( .A(gray_scale_2[6]), .B(gray_scale_2_s[6]), .S(n30452), .O(
        n13567) );
  MUX2S U32829 ( .A(gray_scale_2[0]), .B(gray_scale_2_s[0]), .S(n30452), .O(
        n13566) );
  MUX2S U32830 ( .A(gray_scale_2[1]), .B(gray_scale_2_s[1]), .S(n30452), .O(
        n13565) );
  MUX2S U32831 ( .A(gray_scale_2[2]), .B(gray_scale_2_s[2]), .S(n30452), .O(
        n13564) );
  MUX2S U32832 ( .A(gray_scale_2[3]), .B(gray_scale_2_s[3]), .S(n30452), .O(
        n13563) );
  MUX2S U32833 ( .A(gray_scale_2[4]), .B(gray_scale_2_s[4]), .S(n30452), .O(
        n13562) );
  MUX2S U32834 ( .A(gray_scale_2[5]), .B(gray_scale_2_s[5]), .S(n30452), .O(
        n13561) );
endmodule


/**************************************************************************/
// Copyright (c) 2024, OASIS Lab
// MODULE: PATTERN
// FILE NAME: PATTERN.v
// VERSRION: 1.0
// DATE: August 15, 2024
// AUTHOR: Yu-Hsuan Hsu, NYCU IEE
// DESCRIPTION: ICLAB2024FALL / LAB3 / PATTERN
// MODIFICATION HISTORY:
// Date                 Description
// 
/**************************************************************************/

`ifdef RTL
    `define CYCLE_TIME 40
`endif
`ifdef GATE
    `define CYCLE_TIME 40
`endif
`ifdef POST
    `define CYCLE_TIME 40
`endif

module PATTERN
`protected
]A[2U;R(6fM]A7U)P<J[K<&]^MG1e)ef8M#>X1HZO,^Z]FZ,e3+E&)&7B+>YZ\SZ
K7(3CJWAFM[7,M,<0I@J-RG1]V&eNT^O&g>23FOY]BNJID[W<X[AXY+\DYg+.NN9
KDP>E)5f3N?7_99\7SCM+KCSE0d466E^D<8c2Z[6SRSS-M^]Z\LI]<D)5[b&8F/Y
[X.Pd966(L<E&.5AU[&N2=W,U\Wac^/<))Wc:NC)38<S3,f]L_1BXKd=MC0F6gHf
G2NV^,QGHSWVEBO[\@I[15://\L)G5-ER@PHMV@S,(RWO90(Md&)WS>b,NBa)\>H
XIKQY500MF:5dF7P[-@FSEL,+M_K+CAI^9Uc/GJCaC#B88/(:]L+X+aO(^+8HFQI
J.STZJbb+XZKdCaDeU65Y_<&0\:CH.b4COG[M-8de5MJgN)^BSP#c#PfCX^a9b/7
W./@^\;(Q;>,/JW6J,b[+1fG]S\??L#EN@99a:Yf@&:>/Z9)IM^_(J\G=#D?&A+/
.7J7.BVIc+RcN[cHK_PRbF<DZ<15_;M?9@J(GCH[QJU?1?@T\R1(#?<A]5I0X+44
&dZIK:SH]CJc21^0a.0MS?.UC6JKC.2M>..JOE)_Q2^.A>;-18=--?;&8,:^Pbg@
M1bZ2T-+Y7U?+YQ<.bEBAM2Q-]SggQ61@RaO/g;;cgVP1:g#7\7e)U;51G6#N@AQ
,.Cd;1g.@>94D-?cb7f26g_YT[2LG]Z70#;]:C>XP@e5EEU27/U>.-g=YF01ZS((
Q)B2)bF1O0EdZKM_FNUNL0.g^d.]TLH:O3T)15:WQ.IXMW>NZCTHU_-Q3ZEeHBdZ
]TMKDXM5g-cS>1)<GFG\+[YESE\gY^>8W?ND0fg0CPB_O(9ZM#O?WX2E)O\+Z=MD
8_=@Z73b]RU(D>MUPc)83V8_/2Z@L:#L4cC1X;Vc;=69?C4;&U^+=7+SZcB&IL9C
/\VaLQLQcW6^#g9]@#L4]P)92^T2b8QR8KF=IAYS;@@K4WU9@4[K\1ga;1IJQ?4e
LSaO:.a[RBf\BU@W\DQC#Y0fB6.R,D61bRYc+e5Nb/7TX+F:W;Yd0T?GD1;NBAD/
SN4SWA(M^^4\\gg=&f)-W=:I[+\AT-,V@T]F;>A:D^.5UDZ&Q&N-JND:HCM;24/f
D<OW0M>J-NXfT2+JHdG?8NCQeCI6Q7G9H3-SP+2K^^Dg7:+QX5(.g;BK>+/H,bYZ
=K,EdQ8RZ::5RAIB0U1:dE--eO24V9W[;3I@T?>N?H9M1\,KUNU&]UISd[b^VPN7
4P;IPEVKS@ITXg/O8C#B3WdgB7\?#?HB>F=5,b@D7U?.1.fSgOJ\YD0^9I^AE(bf
J9-_GN)NV/1AV9C)VJSe:BI^-a(SK<d\Gd10Z_V7J1FBGeE^AH[Z10,:RP?_9e0(
Hfa.E19Tc#O,7UM&&V(4V91XO<C3_ZTe]+5S4[dAK5DL^1\SUbW>90GRHe5g[86\
Z7@ZFLUc^]fDUUbgME67^+#K9eEB-c]e9#TaW5JX3PU,Sa_>;[<D=<)TMGY&^O,W
c6Q[+Q?IGa>fF+Gb#Za\S?N(ZEO>X(<KUX<PTC.6a>C<c706eYQ,K<ZfgH[?AVMT
IW5UGT,D06)ICc#[V+KZU[G78:BQST0S4dWb^=9O#b4PE:]fJPZg,8)Qa=S)eU4]
]SU8dcLe6+3<3CQ1)\U6Zg9;G,9ACTLWJa5(N[:cU]V1)5>=88G2QP7Ha,\J[3.6
B\GM]bc5fD/Ue57ZdUbBD]O]?C)V)Z-CbY(^-NWWR-Rdf_eRaZX)O;;aaf&3YG-H
RaW\)gZEL&94X(b<L:)-bU:Y,O=FKG_PI-O,H/,4M=Z8IN5;#T\IT)AO=:_gEH6B
5fU?#C^KAL4>4?JXBH;@>&1S8N]Q&eX0?S[@3OOX&&X(a(-9TW#9UPcN6Ha;bRV,
T4BDgY5CbBdXZa?<4NT-PXdFKEYDN=.-8G>,7Gc5:fQ+IGME9a5RZQBF3)g<-9VB
>d0S-_)@EOVZgEc6(]RFR=+,A)/I;<1OKZG>S3P8[=V2Bg@[A+LMb;<\SYWe\f,9
=9BNZEMNR;ADKY/6RRS.0]DJKa&.P0MEJ2/JNBG;^V;./[=<6P4L-)#210=+\C\9
0Pfa=X.J3#gJ[Y&[bBNY#U@a2FC8A0>F^C,ccD.)0P?7OZCPH3_.Z^B=Y>a[A(1R
JQ;ZDYH-?H[7OIA&[DGad7O,59AU>\egP:5W[DBOb+YZ_6;2>.EX<)M_6KGTdI_F
g>[#c@+Xf\PR:ZcbV\caCH)<,ZQV1:T]:CgEZWCDFNT\7NCe#UKbDD8Kfd)>0SUP
\+>Uc@:PAX8.49FM@A(c7@F=?VS7JPGE5SffV^TK,N&Ha8-=f[&5&9O9/e0:D7b1
?D3XEXIZIT1fWfZN.)]#/^?/TcEI>aOGN\@UIR-U0?WXMZ4&eI\9P+2_90=PF]Xc
4.IR_8?YAWcD;?2R(44-\_Q\4#:)?bEUSI<>bHcXgKKHK+f]F>6KTfb&?2S.US=H
,-;R+M^QbAOEN_/0(Aa4-,08S)1]^Y@JM#,Z/LaY44WD=NCK.X->b&J,)1\\4P=.
PG?9ZP[-SVO#RZSNPg=:3ZVa/KXCCQSOS#gg5Ped9JH-6_\.(SHFBJ\O_:R-VU..
.30TS;(2Y.>5TCH/EO#fWe<F94[&JUQIQ/a)V;FF]#Q#fNE<;Q,-(KJS+:KX^5(>
O;>?79MXZ]C:NQM(C0[ee[BJ8e-[V<,E\V5GG5f8B-4^E6>G--c7fD3gZVN20QCQ
(W<AVK:L(Q?d[V\K5<J7P6&^XW1:IV(NY=>@OeFFH0ORE1?2]E)436J<6bcdgB@e
929MEbZ8-+WOe+A33/WJYJZ+bO?8V9JQH6<H_H40Q7g_5[YZPVb?311\RB,IVFK2
Ob)bOBW=F\9<c/]=T9/6U3c_B6^R#QdG<1UHX<A_Qf.52P;-M.\MM-cR--g]2O];
C/MS?&D\Y5;SUY[U4;b,3#bbfP5)-35MVH;R\XAB_d>;7Yb+UQ:G^HNW?-30^Y>N
5afT+_LG3XO(KY;)A9GE-dYH1dY..CI9DAG(LCWL3JY#2Ia1c0X<O><NLJ&@<b@_
P#+#2>5;>^bg8?QM)DQQGP)+[Ig.8dd/#V3:,eGR20]g7c&O8WX_+C^BZV^]1f0\
WV)&]MDT-caa0DaSWN#fIaP_7]@.eUM=6.[NUaI=+A,\(?9EegF1eJ[F;4dW3^.F
WGQ],2O_=7Y)?LTU=,1(a<C2GJ&KL0IEA2A_(XM94=BN^eO@SDJUe2WH(/^(.EML
(C#;Q@:):((>6,&IGS..OY2SgDV)EHG5HM^3A2EG@=WUa-(X^b<J9dN^MRR.#^^9
AL[c<LYg7W/2fWTB&9T1R?4,1K/>U[SC7(cZ:#3N#8WXJ\d<,]INX]K](g9<G^VM
b5XC9R((C.R/&[)456ZD;8L[^;K<=\LB;#cH.K-.Sff]),6?[-SbT2d_;\B/9YR-
7SI-dg7?dP+:6-J]>RcVaF].(YZQZ@b07G@#-+a[QXeF3S\D]EUdIc\<.>g^)DGc
K[YCfR_7+XN-47JDCRPLGd,BgZNBXe.)R3FC36CE)<#O-I2U@??.<MVO<Z^[a,SB
XeL?Y[08ZX;4OO)@d2b-abT&FLFR&,C-7_O+&DNeC1UfNaX,b#?1X/]bMeIAQ4&Q
?PKCH69^-Q(DG>(UBeGFdQT?NJcg;Qc<AX^gS)d;FQS1gY9e-=0HeGRf,W[)Y0T^
_7Q3Z424=)d\Je;N5(AYBcN4Ya(R/N\0+N4;A6eHdC1IW62B7Na_KH;K\GgIYg4V
7H]g)V,UM8aSG)QWC^[,R>DL9MQ?<D+Yb>Q=MY0-N#O\/0;SL/U=@BC\d#eVb;X9
<UU@I1P1gF=9eKd&;]]>F(c5_(-H2=4\aR/6G,J@b/8UDI@KN]FM3;VN/YT(R]0e
DQ-ZYK3DeIA6ARQ.)+R(0SUSgC+#R^ESD18;#PYC1Y4X.L+5J.&:8SV,bL;S/K[&
8X\Pb+NW<E9/Jg0.]817;+F^DFQ>K@TDHgG8PPWZ<[(XS9;;\Z&3ARP@GVYVKVP>
4cBe]3(LI)7;)C>f6I;9.)1?EA-1?d0f2^G2TS[W@##L4#L#9]X@.^5P\JbM\,0L
DI7U;Lc.AT[(d3U82=H:E7<R3d>W=7)X68RFK&X7dM6/JdFW9XGLXN=91+I7[=fA
Q<)-+dg8fAVd]aTfEgg^N<Q(:[/83e:WFg(b1_>]+;V9D//9^RN/C#Va[,;)(2JS
XF52=_ET>G.1NFJ,=cFSU<a8>X2Ha7EKAfEQI<T\[TBg<:E>)gO#?fREJ_YZD[.0
?;^HgK6FIJ9S.Z&:/L2J8\FAb142XFc\FY@B(ZdJ,BIc3##P1K=fL@&U-8cg9EI]
?LS)K_)^^g_VXfBE\R-\0561+AI<G9gHK^?3OK[M0dW.)?Jf9KU2-5,2>FQ1XR),
6S1L,)[CFX),6f(5MIF.Cg1428cRPQa36Yc2>BTJ2&4MD.bQ;[\6168Rae,=(MAX
F#FLC_])W87KM#5dLJA54&c>A:UG693_YSKW4gP<=.+(G@8K8K4N]_:<WEL+#?)Z
CYZA5dAaFb=H3_9+O=STHf=]cMLR6.D1,30b4=:.bC[&8?T9[@W)bH0g\^?JbH_8
6+K.8[:HeGD:e:6BNN0&R6WSDc#)M_&+DDe&PTJG,X&#Q),J8YX5YVC4f@NYEaR8
=EA87T?D#<,&D&dOW39PC<ENL&MIY/ea\CL#a<Cb\e7#Fd<U@.R9;#_(GPf[DV3/
]>^#=F+Re6LBad#fE.M(LVCgUR>DUWEI8[W#(SO.MH=\YG7Wb9/SHVR1^^eC=Q,D
ZOe?C9#,WSGU=OdUcRU<#>X\+?d7JTK]OWR,@QG01&E;.>B@9P:7N&^F^.0#GUP.
X:K(X;c5O5GL.DY>g3R_]4Ua]IV+FV36CL/S[P=[7bTY+CVDPfCJO1:S>WFPHAY>
V4#LWSeIA-95Gd91g#^AT+YMK[I:+2H?/_WfbV9D=RJ,C7E1?W&]18g5&DAQ4X(U
-+9XHD7[@V5fR10HQZ8&387Le[DaQU9MeK&;F=(W7;/ZQ4:42_]Ca8FHQD\.<;(e
V:(g[84=gKS32.:R9S@Aa?dN4J3eRRFe)#fL8A98PK:]YC;eMcQ\G_&)23EJ2(8&
Zg5WOPHT@#Md]e]RXeG3^-a#?f]eC-+W0)@EGBQ/ZG]HZ(V&C83Xc1#TWYIaK&\/
OE.Z8LG2dgBF[7MY<CPB(V:;#]<\L+5WBeWWY^RRb[3?G=cVQ^F+R)P8AR0LfY:W
GE1a^,C&D7A0>8bSUH8b]ML.)F2DcXR8K</OZKT//3E=WA9@UCIH,E<(O,4O(_G?
T6DCMLODg(2YG]6&FSg5d<SGFN34(I2ZULP&?[c2P0TgA6XHH7P4>)W6:ge/]>Wf
.Q)X6()dO3EE9F7\PN.=_QAFX64,J-+F5(,P5S2e._e6<eBU5@QM<IgT;=-7OafL
LH=H2d^XbT?(O_f7c#a@I(W9+EGO8b[E?+Q(6HFHU;EP6\#9KO,5RIG7J;<?&RMW
2HV?H8^S+2,<c<1VfDFIASPS_753AUN<2=<8ReGRU84]QO--1-.d=5M^6((dCOa/
I6HcaRM+)(^AV+T\OEZG<5d5F)_A@2U[_SVFZH:1S_VacLXSF,&I_1CL5E4A>31.
,\_MM99gPY\ZP5g:)aJ&[,;d43:VJXBR)9<A<#L2^AEVcJbNZ5U6RC]bS9-03T5,
e:Q/:GXOAZ6W],]6+ZfPcQ\=>LT0D2g1>5e?(#FeT3Da?Q+d_?9#_7S,=bfd8d,K
OeU:2T=HD4#@74aM(2O/,=(L<4R_a5A[1OI3:-VWb5XB;(89YR5e8Q58MgQ8/1#a
<eNd58&LD<DS2+RPR15dJ,+Y#[S]<Q4_\^b<N65B[6=aJ(#E6B&Ff#P4=H)c@Tb3
>ce\S(:\4L.W>f(&IdSf0VVMGBRW(0GUN)K^H@=F&d5=d[c?FdU<,E\M2S4Y_=6K
+(;H?<)W.1(1VURV=VHG\B7LJT3dD460CW/@+>)Rb\^_5F9C3MO-;;&AXda.7bPE
cTc)A<<fGcfS5E0&-)S>A(\;DTNH)SgZ(Y3Kf0I(5B7/T#-.]M@.81:RDdE1MF3K
3Y=X6Q3NBIF6VCQN.X6d?aP5-<.EJ1T08MDT,?;42P@JO#-\P6D3<<.?)D1,SWbJ
315PY-IV^C6J+4GSU;RVF=^>MbL.(E)7Ye/TU(+&OEf/EDI#M9;2#+e_a.Y:D=(H
4J;f8Za\2Fg=KXF.0[E+=7M4#<G1(B#9)&Qe&.T],59,(IVfH=)/]eZL9>U>f9f(
UFO[FI:ULHd0P;a;H,-<P;=05^e9DLM7Fca2+X-<C1PZ?_KA>6A\3P-\EAGG3T\F
^5b<_P-6eTG/5T(Q4>b9dPf?-f/OZF1L,@0+abdO-LDbFN?U=IF&[3/677^ZfQ&O
-JEUY)52L_CF7e[cK/g<H>BEND[OQE3?:GE^T#;O@/K)MIMNJ6F\Jc#f541,O3>F
7d72HI5ZAOGQAUH,3:WbA[O[1&c;3=<^,HSILJ+]=WQb>WRI5=T(W-^V:dU6,H@9
CGAXA@^;/L)[LK<Y4a#V&+0]>+N0TD?.^]FCE7:0cMTB[KFHNBRV@V/WLcP]@c0g
e4[HS(=>e^DZ7#a5U[G4-]eCKDN/Wa4XKAaD5I>ZW=)UPE/FA<0R25DT,59J(.gU
3,0H]Ke?TZg\OHNVDBZERAdXL6CI)gNC[-(/Fg>@0BYE05IdFG_YN#@fOV\00N[?
:C8^2AC,Y84#WC]8L;LaIK4f5Gd=bP5\F.;FF;0.Hge?K,]^S6;U3UI5&PSY)]8U
VZ.RC(V=2#^bYHb=2>#/);,==.7/DcULU(WV>g#cCPf@<L#E\aZ6:cB6B[e)FNH@
X@95:VDbVN0L+_TQC@VIdQbSF:S1Wg1HEKd,81(#-PER9b04@/&VMM]F1M^Z#6B&
K/8D-P1UMb3?@RV=ZMagVER&54;SYJ;Nd4L=FDNGG[KF)7,3e4eVP\/dNHNE5\H.
KPddL9;e:DBKD&ARCF(3MF@)[B63Y#&dbdAC.QbY97TA8gN:gHR0H.aVOQ^Z3^Q]
f)^6+ZG;I/H=&dBL#+2-4YXDQ;2Gd2609P;G5Q.4@2E.E[,@)A^7f&VB>2E?:JGW
AB4QbQN-+C7=5E5>E(K90B(f&#GXZ\0B\Qe,,J&)>6d#WOHPC7W4VOD28)^@cI<Z
RKYL#48]U?L4#<H9(R@._5g7FCcC8-Fe&@?/8T(A^Q/9K&E>9IML-,TUg;&&^TD?
=RdSHZF,-\):aGAWR.c]Cb)gV<>OVBXX:<KdEAIeVKSUG&N_#X[-+(NLI)DZQ.J3
P],S7ASg5-[>Y800+eQ_gg16(APEcC0aF+KD?E]0>#WO8>,Ib9aAe6YV\>7A?5DE
8g#]C9-(.Z29^=\^6B6L7:&HWA&M(D7E\HUK.#,bXLQ36\Ed>ac^:+0@S#48<6AO
JO1IPJ6bG0:\;3[M<Q<)L?-H/IUL;7Y;Fb9NPd<6c(?E#]>N^5(=Bae9M/U^c:G0
<R:N265YGM\[J>e(bO(#:EFXKcCeG4_R/R:cBS6G^V)b>9+:+QV[d.fOe-1?KP,/
=ed4X<[,B67/9<eYTE4@>G/X]L.KO<4Mg.YZ>S0beFXeFEB^-Y/UTY)PL6-;4-Qe
b03&=RC-^aFBO5(61,2]>CP?EZ49cJ3G#>#AZ#[Ye1:=2GRQ6d?a,Hea6-C[=I1J
^4-S_:ZSWY)G8S8CaaK<KYBH_-K1VLFSBAD\^Y&YE1f8//,7\+_XJ^4K83>G@)ea
;,g4a+[PQ=M>P0(I0+A;b25URN@D]B1e&Ja)YRY\a=,?@D=XCS8_F4T0-R)GKXdI
>YJf?AHWU\9eL<XKSFL?LD=68G?4TV4RF?;dAbNE2ObI]PDa,gQ09O##Y=BYZP?B
P.?;,)?=24-\&(<UB;B<,I@R0L;5,.Bba2HSBI:Z7P=[;O>_FDILTg9+O5D@BB,b
N1;e7N_1,d/J^=U3QP4T@FFeR0d3&AM3P[OdTb@+Q<2K32N@9-HV[B_\5\[\V+K+
J=;@+GcMQJZ4V<;QYV]G]VeUg7M]f@U7e9\ZS#VQ.A)IE./Vg8DI.TZG]RgF,OL-
PIX13P-;#f1#:V0LGU&W/T3?M5B9Y.FR2N4gYU3WX;].E=ZZY[E1,;H4O7ZU^FD^
d5F&PCUMYWHfPGI^g]H[,AD^18RUA5(0bV:HIX+#(e&+T(DV[dSbVbeUNDc976>Z
LFbgB2D54^LbP&F255S\@c=@=.PK9@#23g\aF1_d;A29ZV9H-&6+-F=@9DEU;JaI
GHH.4;5S(Xd)QeRb:Ia1DE<Kd#=HB=<,)XV1R-_)29LK7^e0&:JZY1\ZCb5WcWfB
GCa^WMKWb:^KY-RC2JNeg;8gHAVHbQ1bOH+6X&E?]&<0@TWKEX.2]YA8c5PN#3c8
_M.(PJ&]SLfY/bQOB@^-NWgPQFgPNX2I);V>B_V[cFCI@1CC1\6U0dWd09=Eg>U2
47[;(<cCJ)_d(>A?f3b\AKFK;8];D)&XfKJc8\BbK3)AWE_JECZ1+:MPFI1X<5:P
7c\Y>e4107NY_:=c-_c^U-Tf@O(Y;R30(WH>H22R8Zg11:Z04M^.L>B-V\BAL]/:
S+TM<6O6KQE62]M.0VEB2E#2^I280X:>-]4V1HOJVLS9=aVB-:b>#<fVKMW-UA]_
J/S.B/_7LI//8>A9[/S:.M)7<U>OTT.b(.+=JB[41W/5JG7ZRaM4aJ;(:ec9@I3S
\Y^Q2,._>+@NSJY6I1ZI7VH#L,#ZG>9=c&TL1g@C3S=U7<G:FNd7BUWK,CcQK-b]
E/8SI,\16-;0@Y1a781X45H4HE3R0&ZLCA2LU(b<1<]H=2_:gF=^A.&S9/W@(;]?
d(d^941(].&/6(__]ZGGO4H8J5,_:CT-?A1-CbD:8G__=TQ@4U#PPZ(GSNC&J8S+
BF(-3KF5R)AG71ON=^4&+g3[<7M8SS]HUJgAc9?WZ8#5]JHW^99^7=,fScSeW3Se
3[X?bXa8.?aM#Y3Y@&)_B1(gJH];@](f<_@N&#\cZQfV)7(&Z&W41JdA92,DU^W4
K3^:&R#\Ib)7d.bgWDG.5c=4AZ[)ZJ)?I7L?P9U\E.P@&\dJL8<e=V>40/M;f&0-
eH[[S_7H0GMbZ]8<:\)fNZV=>H?bBO^.<dgFI+LKD.+<),3caeVWDLQO91@23E4?
<TD(IT>FgCe&.DEQJJ#-c6g5=8^5SRX2MS>bMTRU)M:UDJ-I_P6U(Mfb:2<23f-U
dC:>D;c)N/G_-XXU^M-KKXLBK./QXPZ;TH<X)9O5>O-)^@-PY9XaZX@2F?@<POP=
6KG2DeX)1.),I]A^V7S4;@J4fL-Y?Z/YMT91K/aRG5F9FRcL.\TaXLAJ-?@NNB-,
7g0JN8GY;:\JA?)1a]#=YBd19^R.Yc<1&^+E+U+NG[)BNVOOU1+/,K8Y3D72K;a_
\Ef]N7_(D[0Sa<aS>/^7.W/E0)+L>bZ7d:6P[CI&Q9(+Nc=bY?:^3&<A?(?#0f0O
g#<&H=PD@<8T/Q^72?)Qa8_e#HLTN^<C>G/3S];?N@V4OV/:@B+b:HU>Z,GP73W,
J[LAab2GP98JaJ4D]@bEWAUeUJKP+&[I\HU9N:\;1b>(N-JE,3f:I7g)]NVa_V/J
&(:Pe]/FdbWP3289(cMcJC#:3Q[U#C8SL+(eM&9GMZH[e[,5-I\3\^H1b2L&fMJZ
[Bd55]e\&?EUW;Mc,FN32c3^X9D><#9e59]f@BQABB=6VZUMJNE/e)N6QTH5K.P[
1\Vbe3eTe]/CdBF&<c;CY_YHGBY23]g>;_MGJM@M8H@)af\ZLKZM#ZF1#]B4M5(P
LFPdGJ-cg\Ra^01(bGNQ2\&5D=+5)M(#C;dRfHB,[6,:+R?_b=]6\C=:3K1Z&Ga0
e<&T.9I:W>O/O?eG4C656_9/:(eE3Q9>>9;SOg41S[5>:bL8C7X8&DL/:22<@M\X
gQPLY<B^bIKa;PTN5,=K\J5=0-bIH9J:?1(D>gR8&B@eYF:]?C(eZJD^f0L3?bP&
eV.<_O^b#MSTN#IQQN(S1GCYUSZa3f7@@Pa<N^U#eAQP00I\I__@J334:>4\8VHD
2R?@ZS]af(Fg?^F^-bJHcC:.P:^K=:]=)A4H8J9YD/NQ=0c&gK=)X)2@f0_/dWS=
\&&G1Xa]FEU>3:R2^S\D8W@fE?M86)a/\V5>Q.d?3E3Vdb:XcD[>1^fP6_FCOAC.
D48Ca[X^S\)BPZ(9eP6NF6RbX@LM=F+4N^BHO#>WV#@B(\7_M=Z/:GHY78UI0D.O
<1XDC;Fc-@7#Ed<a/YSICO55N=bR@9I)X>G/+M@YOeDfd-FPU4;0C<XXH/JddXZ]
d+V=8c&.a#R8TW3:.M]AY08KE8I5Yg>Ve9<)A1\@bdS+cfb2V,C:X4Q1RX30Y>5L
1\FC3\cUJUC_GXM/cQ7&7Eg.FYdeYVR=)354\MH.dCD:a(0RQ-?5SI,4M_DNWXH1
=OcLeQM89eeS4<2:W5H=1K;]FN2^5e2C].\<[;IW(SV9HV5J<^;cL#?#C2P&:?E=
W(C:6de-CfJR;9V8W@7ANA6+f@/_?).G.\\Q6G^Ub8ZYJ-AJKSKE8[Y_Hf33KO.5
<UP_)c4]ge,_O_6WL6>]0(V3CaM=QM0@I9?+KbeWP3\\c4bX&X6YO,Z#-C0Z4eIV
+GVT+B@N?H?-KX4O@:?W>XGfQVXS0D(c@I1<+E]Y4J@)_VaC1G1G8QUO9L^24^PY
YK>\>&b#(2MeK1-TdYDMPg1d(NYLH=RU/f[+-#Ba9ADd(=B]e8RGa]&eQc04?Hg;
\&EC]Q)XY&aLX(V4[++L;(.(8Dg=/ET/fQ\e1LLO47c0_FNeI6Ab<Ld@0_4OWL]1
1f>;M?S1G/&NZVJg6\dWY<Jg5U\R/aKe2Lc@)2P.g>L70IbRR6e#C]=3,^feZZ1D
<c@&>b#+LRNMA6J6dUMAe#A6[CW4IV]YPGfO1,ZcOb8)@+[/)d@GT7-?LeV1(BfM
M(,M-QLXfXQZaPU2/3,2<fEa2Ga&.^)Obg@Cd0KRXB0<2P5K(]\AQA?R<b991S@-
47#TOc4c6446S:OdcgM.+A=#ZcT<_da=Q?F(EDEV\]::3f+aeN?BI\RA(I.85I:^
:[9[b3Q37+B#f7?f5#Wf&<(\@gP1(O-<7X_+D^;<VL];?]+AK2/fe.^La5EP:R7Y
>2[/VK_32;9#eGDaV.)&_[fdL,]K7MFT8_9#4F7\N7=PSIcO^:9+C_&a4Y1+eS=8
\NF,:Q&;=agb_):Z-#ME+R\BP9(g.[bTd?G(.18gP;\K[]9PYQ<aEZ5c?_a2JH<#
aedP?2K=V(b]E_d(S(()6ceWafN;7Q3[2H:YW4J7EKH)PE6BbdH<1UE89e3P558I
WYc=MUL]6Y:>:_BI<.O7<8[U,FVSQTB&Xg8.gSY)f:HEH/Y?]X+F95-_/\/b=3M0
XZ?:)IVK=NYe5&[Ob(C4Jf#.[G#3TL.O1JaW;U2Xa]4Ya0)R&+45;E+>/D8Y9=TD
,(HC+(&DTAZT[.Y?EWRA(3=^=CU9\#:O0T48fGZ1a>N2DF;O/Ma>?;d7@NO-V\^0
.QM-)cX@29aL8GIIB@5RJ,eF<K//^/aCR7D/YB8)@fgACd-FT@:_RW:PG9E9X^c=
3E,#^P/c(23#AN4JXKU+B#8Qe##_cO6=];]6b@:&,dQFY@4RdOGF^TFMJ?R#/;F9
OE2_J)TaN5Q@Z.Na?VI21A^S>O_-W(LV+JFJ##Lf770a)^Ye1,UCQLc\1[G#QJ+G
?L?bQ2:)ZC^JK86eDZ?&&Bf&OW,R8G7M5Ba6MDCKfgK,)_(N7]?)I_N\b1CWYNHU
T\2;dJ<3Y7L(1F6:3C:_A2NXL#,,=CKgA,&<(cQ&<P.4=BC7C=E<;OL)XZ9-.e;K
65Z3<;T4T6_-YM.WYbUMQR<7VXPICYOP8P/ZA9Y#X&bQb:0O;FIZ3@/P(J=H6V\g
cF9N-UK3VNg<)[K[N7:/T1R\I=:40BIKFBV[/&E3X@cVZEKN8dQ?A358TWQC2LP5
-,0R96EgM6V]a)#&5RSE^6fNDUS87BQ2fLLL(#P(fW_C65dLT^?#aOSXN_4=F=g:
N:[<Oc?e;\Q1?GL+KZecY=dP\.B:D?5-+E5D)PGKI]1F(5?bCBQAMeV9OP9#@YdE
,aP:)V3RHWH@MH#^/@F_MIIZF0G>\HF;.HdfB4:B.5HE11[?g&99S.;PEB\7(aVJ
Uc-;^6C9B&,<1HOI8Z?3)4aab>NVSXRA\DQ,7JbAIS0>VZL77eSM0W,H-#@#2\5g
=CUQ6K+-+dLO5PO4<V[KZ\A#fXJ-Uc&9CKJ[N;FA5.>1SdfJGTH]dP2:--;59B_1
^/NG;&Wbb7>5-+=-M=US5N,H2R^aDCX;>F1<>4f(aRRQBVc&&P\J-Sf#F.^,Q4f;
XLd@2c3dCU;]]Ae8@[Z^F4N)/9c?.H#_1@?I-M,)BR<3eN>.#?YRea]Y,b=Ue5>(
YaF?a3:dGLNdQ>>LU:6Y3-CN_c9#Z>)X=#(TXG,3EUB9PJGB\f,(]G7,-(.G^SX>
dd(4<E=J(<_fQI,HII,7(CQQ:P^HGF(?f>7OI:DZNce.[)gb<aB#9Y3JP^D[+6e>
dbd3R=W__=_T2[=-2LZWJ/e8L(,PJM?X-NBK<JX>FZ1\2.H=41+0NI(g,0T]8dG?
_]U2aVI;69]AB72PP&g&>SR.UQe2WPd)fR:<aa@CH9W=/PIHb7cF[TRAI+3dg7SP
OS_6+Eg3fCL.:_W3SXQMU_WYNM,NH+?9X7)/#OX8D2HJH(@UfX8:CWH\4YGV:]J^
ce@K>MX>&/U13;0S<E7>=/1G8ZfQ;3c16-:-#_JCJA(R]@gcU9QE>Z+FgOgQ/XX&
L?U3;T]KY(98f.,VD,.LHIb_KJ^^6<[OX&):JBOASc>,67Z6[LGQ8/JcT[R#D=2(
5a;IE4))_#=3:MHFZb:6E;BYW[bFS+\7[S5<g<3^P/WcWd[=061,=;@=/V2g;c;M
QQSLW?YUc8>>6Q2[XYdMT,:O&BOW-PZ_?YdO3AC3(\d9LQ4RFTe&bbQW#gP<H(U=
8:gN;+Q\H)CIZ7b77FMC1W&]?A^96R@f/g[1@K),NCEH?Ea=7TDEU^g@Og4^>@@a
H<<gN(FI:R8)fAggKVG)Q6U6J3.[,.b?#,?)UO1c[/L#J@2^J0X9=@7HKDAU@BdC
<K<5B<,.f8B24VT,KQ79=3gW\P\J9K:IFdQ_KbgX\Td,\V4EbEYFd_I&Qa1+fgM:
VF(<3JC4H2(aeL+Hg7bKf.7]c^Ld)C#.bBbI6)Kd]<SSR9f>=8GQb?CMG1+2a2B)
GXB;NLUG&^fBMa4P(&FQ+]W=Cb<#PJMfT6X9?Z@UQZ)#]c<))BXA\7@,GJ9Q;W@g
9AG&;/1YLZ[eIO;cIDfeQ3Y?)HF7Y_/f0M54e@_a9^5=39.OE+O]9HXHb=])1:_?
WIPL^(KIFE?.;STI,f@@KPU.[6GU7_bL^PI;DW?Z08),V^#06>3Y[U]LUUKS&fcC
f7b;#-g;WB6.+_5O5=E_@:2a=02\Z)SWRd=5\4?cS.VVS_^IgK>f&+0B2RKQ,&1F
>ff1O+fJR9(]3KEb/\M31KM@VU,DZVQ;YVY\SYcUYd^:>SUR_EO+RZ)8OBUK:H?b
M)ZYK2L)Cc[5^\/H,CdA\DA>M1G@S#B:3Y5Vb1Bdc.CY)12&BS-XW94;g_2^P(Aa
/cdXQ=8F4EQ[LL&B_?Ee#<#;6WMBb@gd6R1c#A#/L^3b6Qg[fY[e]&VaM;7-YA@-
J^UcLCAY=\UVR;H64&ba73NB4+D&CN^X\2XL@PKEF]-Q&@gMCa?gJLT.Wd<1GPaE
BD/4IfaRQeeDTS7gE-?gB3#7T.RTgQ#-g94T[ce2@b54LQ#OZYH/A)H@+;dO-IfD
c@#)ZCfKX8W:Va/0S9fe8JNaU8I;:1@e@.]bSYW4&^]1^HT<40#V0U[V.TY9GOWT
Rg;aS9^d+#f#.EH@M@NONSB4[0.E2<aZbB>O7R#AZ==3PI<M3bScFX,)ZB)[dRC@
f=,E\82W4XB-Vcg[70:QUg7Qd7Q.VWY,((NFa=1dNF1Y2X/]d=&-NK9?L8]R095T
3S][G4^=OT\^]\7-Tg/\Q6@Ya;/6PK_V8W.KHUI<@Mg4Z7BHX>N02PSW:BB-77a.
QR@_]VPYa=fd&NDLN]Sg9VaYZb;J9_K2W=AK3,?f8;GK@SL.3QFfKN<5L4HQ.EM-
O:=P+NXAIL@5[30W#NIGOf>6[b7&[T@ReeQVAI4+Z,H:caB/S:2LfNL>>JU_M]?W
Y85/]^R)fE3/ZFbCO8E<3FLDD4H3319S<8;?4VYS/CIQ>fO@VT8:HgfObA_^>UDE
S3f:HA2OZ6->K+Q6<b][TX)3.4@;QN;?+(0K4@eF@4e#6I09K:\PLTF[+F)L9\d_
A].2fR-(f9-&>X#&LdYd,dO/@6JgY:4MS(/a]g>f,2D=Zb=,-B@SD@cWN_3+[N23
DXO\83#/A\@XH9e#G&C>Uc6O0XF4_6&E4AATBOdO)\;.aZ(RN:T_K0SAV(>WP)_;
^#):_AMeaL@B/(306:W4F)V60c910X[U-VP:eE6c<K_DPa=7?.e[bF:dA1?YOAJ[
d;_)5#@D-N/EN2c@A9WR3YSI]<gAS1F&5CWPHaL9/#:BW[cNS<<:UP<;8.<)0324
ZAg)U36<>c\KLF9HdD]ac+>2ORgL#I#2)U.?&^eUKdXP>Z)7\WWTVbL-&T]=1EW6
:5@O_E=ePGGfXBNYMTGL.5gda1N1-7fR@,_^4T]R.2VK5JKHP0M@#FM^P>&LG06)
DP3A:@0[NdI78Ec6?Uf^#<ADWTcW)5[1E[PPLKI)gJ0GBI2^#3X5DfBFSf3b^e[g
Y00B?S?(/WNXagUY\,=2/LY0.:(57^g@:>fSG-;,^SSAZ<5A<RX=;LKb94^/<NNL
U5KKO2+\=,e\9XH+(,?V1;,X+;ZT5#_87Rce/UgXe1ZPe4Q5>[+0V)>b)D@\TGD/
E[R+7bVEF[[;KWD/(Y(XY2c24Z/OecT(L7VS(LJ-4<e-0aI<AK8g[=4_ZZ7N3-J_
,?f>aE)/.Uf_@:UH(J40fL3\IL&[N/#><(DP8aH,IRSAe+ARP]8-QWB::1577>([
YdK+Dcd6ac+#]FSSS:#11[Q>Q]gg5e@TfX#O]e)16@^66>ZD/8OQfV=V)cO\<NX+
Q[HM<g.gf5YSJ@<MVRVE,(8\g)4)4ALgB#6644dPe#_]B,YH:5RU)QI&>T\UB^5?
17((],TYE&#g>)4P;K=ZQUb6U>Z<[P/dL]=M[N,CVgZ5:(]&[FLZUdF9=d5)eF5/
3U-<&>f>?(XZLNc3^ZMOWWcJL?-4U<#S9Cc&,#+N7<?Qg--//FdgWV(?U2HRde6@
.SDLT2D)bL\H(d)I=.X1L9BX&TU<J5@+Ug889XRfG-9>FRbX6KB&1G4cW\F5=4#d
3=8c7U=[;0aII6D@01I,c>]]Sf__c<HK<c?9E?b<V/+NQHP@e7D1+P(MAJa1WG>@
c3>Zfe_#[](?VBdJ.BcaK?d)#cXg<SOaZbLb9[4:ICT>_4E2-<)fG4,-^aa:fd1b
&.>g,MfKHW#cDCZBNMdaIEHFP6Q.5MWY&7O.1JIgS+ZV6ZNO_a[DT^?RTJcBU+)0
@LN+II<TXfdTT(#O\F/C\[DfTf]C\(JgV;I&@Z+,>NRTPLU0??52K4UAMWCE/JJ,
ER3_d->H,+A&:#N^LVfWQb7H3TR8P5f0AFAFLM>IOC25?@\^J/FJ5Peb13VF5D4D
R0(4)S^L7e)T,:bc#85cfPO-11A=b286HL.^UD\a8L=Fa<2:?cR:&<\#OLY4;fG/
-/,YSccRWE_LY1Ya<(Z^Pg+4#J5ZCONBEd(Be+D9+e(XT_^\::BRZ@6;#U(I=NQ:
A#f+8b56DDR@18?,-bA2_]\HJ0JHC<b9aPS2:LLKMDC_#>;ODH)beLW#5c;gD]VH
VRQf)HaRY^f4CQ;d/J@QPT9@?6,D7GIfdbLR3#gDWH5a:_,cSOW7RY2[aJTDC49c
_eg@fFa#QgfZRO)+CD/88#f+64OCV=UXNfI-5KO/>Y>GdW.9VFaQ,]D0,9g?0^3c
7+A_.>[=G<WCRJ;>EO1TPO-;B\[A<]ZQ#J+#F^.&_2C=2GKWe7>\D??,Q[:E];UT
-3ce)WaC=bK+a.S+W8?&gg.\)#EeQR/,UEMYTMd6Q?bfMI=#/VIed>>8M<2S-[/X
PI8PgI9/&WW+L5(IFCF6;P]WA_H(EZN2V#D1O4;7.GK:9_^Bcgg;6_dD2CWDK9<3
V@a64f2PZD+4=]?#e,V.)2^^&[QMZOU969V3SULD])L1)/+VJ8WU>Q::WQ:NE[OU
V=VA[8_S&.#FR9R8/>fNB[2eZ^D;LE4PP;;)YTbAN#Y[6^bYIXfTH(3[>=3B[&;N
E14+2Y]>7c6KJKQZ&OGS<L:GM.N80c5K;B6+4G@K,P)RM>9Ief9:HYQH>bY0<,.D
0D-U?HKO3>T[e@0=X/ag5Ea8gcE20A\fa48f6O,70WHOXEKC1A.d0FBbUCd_Z1-K
V^CC.&LP/,cV6I40;RUHCAF:I9V6=ddA+;;_;+KCHS<P+ZaG[7a(?G(6Cb=N;8&R
:\V>OII=9KW<2<WOHPMgJ@NA<2?S(gV9M=6^,AWV1G0#UT7&S\3/Z_\V15XU)<C]
+W],c^#dEJ&A\W<&A+7RN8E./NEgB3[L@60SXQ69BA#V:&KS@;B?W9U-;[7WDFC7
R@g#(8D;3-#\Tc#gRZ,S9V6P-626:b,Q\H#,E^S#&-2(OcGAgIdZ,CV4:D4L=(YF
ZHP/8AX:aVV803fF:3/@20E7.>cX4+7?->aIYXU6)?)50)V-YFfSId.QK.<6GB?V
^b5c(K^LcO+75U,\,Q;B^:<0=>M=9:e2::R45Le>GAF>N9XYc8SYU7@9J24Fd_AE
DZQRRYXM^V>.<;dU82.KKCKQ-M2ZKY^XW+,7OP(A\QQE,7O<R2N;-?/d^cK<:NRA
UbTZ2@T6IQ)TQ7]<GV_UM9@-_Y.6Wg^:JE880>PPBG0XTbA3F]3aSUO(bQ04c6\B
dGTLXX873ZHDIOE=RWcIf@7Qa(B]>a(]FgQLa@a44Nb.UK^PIS;=+TGM77]KYEYW
PUf>>NCS@<fG:Za3-P#BCaWN->-BBR]NI/:LCI+Ve1<XS:>K<E[\>5&gEY#1JP4Q
aOG5I(dGA\Xb:IEIH6H-A24b>MF9KBO:NN)ES4P]JK&5;QMK)QM.Gb1/L)b]b-Y8
2.HfETd@;\+8NO6AORD29-YK6N@6O8DQS78A</8SO9W22+efJOOEY0c)Y[\IPM(7
0@_FQ;PN\^_86G6<V9cdb=&RC3Q2627;(96#RHT(=R0DPZ5_EA4OAPf5b<75)/5X
U6g:(WVcARQMP#CBP>AdJdT3([fd?+=95^V,bB,72#)IcK+_GX<B9EYgdR>:DS,X
9XdA\2<2E(EAW2f7MN#3[=YD:PBG4^^L]\BGa=TEC_);17^JZBD\9NEFX=[CSF6M
C@/3e4H(_/gRWeQ2dbA>FX6YYAQ.?)R,=ESe4M&Bd6QB:AG=g).=)4(Y[[\20#@+
9M#]GC#P(OXTJ06&;ZD+18YBVeM1HRK:NP?e55f.PJ_8eEZ>a(fC-X,\F(?R/E=6
AgbK@J6U2eV\NMO3+[N0LN60LBS4D#-.K9g5V^@gY)d6)TPR2C3>Ya\+@_E(H6dV
\PV?F@.\?EK<I+/NRC]H?<_-T4/@AGe9\(e1FB8X-D5VLg06V^XZ11I&Nf)ga9Lc
WaNNC<YVLU?<:_JdaaLIYJYH44_O\W[;=DCXX0QRQMJ7ggTg8_Xd]A#K4WZFYXZ<
,BSB=-O0MB/JdLb8&22_0a?Zae=BLZF5Vf;</Z_KNcc8^B3Y-#Vfe4/<59)TCF(>
\Q.Ga^^^ADccIM4)ES]#V\ZZ<>MAYNK,M5E_AB>:3[UHGM40N\71-[;fE-)f/?bR
)SJVZQM?gb)A6+bF1J=C6a6CefBQTDJdXXP@T\K0ePDIT<_+/bHCTg<F^UA(^c6(
\W6SUAcZM,1=f11YFJJbeYc9FPB..)b2/<+O0JZZW7?#,]M.<CPN\Y]c^Zbd/Y,2
_OB=UZS&,=4e<_AQGV\cYOY/+?)MPC]19HF]P>Z(3/WWV:2Cf6f?H=P=ccF^eREY
U3Y8(VJ+UJ&@^66P9/J.cTIBf^.R5aP-Y/:,4(<;4bD<9eR.T_(SP^5/e8.Y6/V(
YC,LDX5JL1g(cUHJZJaGK^PbO.@9_6&[W,VfYD)2?>W2KIb<L1@Gb<b[U2J/&Zdd
9T6Lg3V.aLX#7#89Mc^(4Be?TT/ZY1bYeIDHG8+1ecT:([060@W+LdX#S-CBL/0]
6WcM0-A92UB\[.A&88&2/:0R1SM=6TX^GeT&C;^4IHHQC]:DBUSCO.Qe-=Tg,7_f
T:J^b&e4G]NI5SLS<R[-E.XWMH+R4VQ.D8;@&cDO)Vg7E,cQ1Q.\93LB_@5R4X=#
a6dP(SMRZ3>FIGYcWY@1f=\8YM]c)(M9fKgV7aLYTSF\[DWJ]d:&\HHL3b7M,(,F
_6GPNbLGA=;_;L:H+T#]6bDb7T/GdJ&#6TM/[\cUe]25-5@?60O<25S;0T#b+X2M
TN57PHQ)<Db]FW>PX^6Q8_(V3(X7d41E+;J@5CJeWT11E5(_Q2^4,\c-;J430(/[
H0\&)4_O^VV59(1+11NWFZ\05S/GOc#2^SN#2G4ZbJT&J\82+?\bO)P(0:HJ:73e
W^IE]#@fYDZ?H:&:,f29fUH;[_HAX([M/>QX6c];DcUB#d6)UEcOS@H-:6CTUda0
81dY4F,Bb>SD>UK/@\P;aUgN(MK^3?.@2DKLG8H1,C7EX3HL2/=8KCM_.S5XD_Kd
]Qg&&3Y<D@.dZ@NJWe.PP80CG@Q-)CH_EWa<QQE-,2O#LPb3I4L_2)Z_1b4P<Wac
02eADV70,#\.fE\>2X:96cO^a&_NY1dQWg(g9XI8:?N@,;PF)AU:(TU(&B2a#0;T
A03L=gc<BJ8F;J4aKdeaKb58M.B=e9:GJ,X0O1F\_Q46PAFa&@Q\\2UH7(Fg04\E
YgR&E3O8GFZBRgV2LTBZXe2>aT^H_e?CZ:>N6R2_4bOa);D[f^V7RSMR=8N1M5^&
Z.6\a_1BU&=4b_/E)]?@LC4B3(Q,74;RgW(I4O(#&FA5G8=\A#O.E.8OGVGS&L=8
)JFZO.eSDaX]MLZ7ZEf+2bMJ/U=c)9,dHOdXJXTAK@)aHKeQ5FIQA>:JY4K0gLQe
B\A1?.+;W8=2:=cad@_#:K#9V]QV;5+N33L@#CI.?P&Df:9>+ZE;D7P[GPYe[K;W
;(Z50cSE\_A2NKgRE]/@T#V]#<TX5IfX9gWfO+=2e>b1?^#fe]2E>HcHCFA;0^+H
YLK(PeYMCRQJX\CAYW\E8<aW03>NFF-bHS\O==c[)^H9OYC?/LI#@1<F(L&CV9Y[
G3QFDS_.;:V0aP@4;HEYBeD0f<3;5JeJ4(7fe0?L-FC6&f)CUXH>O6]O,O)a:FS3
=@\^)cSeJ<WK:@5/#^4__2VFg=4<H/F(OFP:/X4R\)]>68#><PHM@NTZ0?Yd9RTB
2.)^3ET3:O<Fg)0M;eIW02KfVT[6N>=R:aNA_ER9,^7TK2PCT>ZL82eWID/T:CN#
C&EA]>@[UK0XLCGG3UG&1Z8aQ.Ad-WYFGY+X(K[B2gRI?N@1aV\VD/((M2@L7F?<
T,OTRU@5E(2(>Q8bWOf4LT6A.QW^gZ5NW[J]N:M:^H0V6]#gZRb3R\<NZ]^.>_YI
G#?ZIbg5HM)VWA0G3Y(_\G2OgEa0R-C?S&@-QcG^@>&cG745FgQ0TZX&Y-9MaTcS
)K&6,XOX;T1=SR6.fbKg-JeMHIBa[B;2S^>cIS:=P8PA(VJB>bUS;W^H<3ZDfO(Q
ZXHDHYF,A^N)8?7YK7WL@44B[XM<::7TE6TQRMd;QXD8?[[@M?S1A#@@85@NA(L&
cPe7d)TXETX8d5.+dfGX>gLdUU0dW]RfJ=->:]R15JDOb.#VcJ]&008#DB,RJGRT
ZI4aP)1fbP<6T]9>^WEV(d6aU8BeVBd=[I28ba\BcEX_)^4-P0QB3WEZZA1>2A_Z
&d0.?3.NKYZFZN=UfR]:c;Y:OCBB\1748d@P3Qfc/ED>7WMB+fcOOHJbN]N5U)<T
?[-BF0H(AW_7gE>Q]P6:DZCQWeQ9YNdJO;Fb3KJ>)g]eA_cQ?U@T^a-;SgZ^6g\;
@,9[M6ZE-8QTXFW?AEQ-C7b1IQAP<L,faR]BSNMXY>)V9J48U6@NPA<LDd=&,Q,[
C[-@FROVAe><]U&.L\&,b1d63I_U87+6.[6MGJ:dbO4;]3@PO>:\;\7FL;&4FA<E
a]Ka9T3^3c@f[&11>J0bKfT9<L(]c@\7EdX/,a@,D6FZ0gbDX/WL,9II^^L7c]J&
<d)VgE>b:N,TSW<<2&YKT@G0Y9UF30HgM[GC8Yb^Q0S.)Td-2(8,J>0]8[42O5CO
40_Z.b@^5&N#>,YE5>e_OHE/cNXXNd@MK&g>3H_Vb^O?9XAP_c?>QF12g?#2cg/L
U4O)LO0#afD6SDN..7AgBGNWR?_8(+B<IF@\SLLFZ&=d_OGVA9;fZdbXQ:L.d]-f
Ia&a]<ECIOd?NSMec3#6>H#+B;78;;KK-R8H(BK)617Ba]_c?X=DU13Z8#[d?>a#
VUad;X[@B+D6#-Pe);IYdUb_19B8V50/4b-KDbAA2c0CD>,N<<PJC\YYL(UU4g[R
.2#IgLUK[8V:HgR>dK0?DH@OVH7RaZ.ELQ.f-ZJ-^(.21W/6)<T&U4>a#&3g(I:-
a/^O&(<;0+2M5QH<WY<U&0MD;b3DFEY6+?;JSHS]E3W.gdRN9R^JE<dE/N-P=FV_
3S^X(P?Kb-1gII[:6dXdXD7^J9#]^S9,/e3-f91GKRZ-c&bAMG:8V?BM7W[/VbT\
SE^,9-?#3N]<U8#Z1K>[>-EP3gYfM]gZBSU;,2eM##=JZX\G:E12N2#N)3(b(BP&
LD,J]]FVF(O9a_Ic-Ze^(H0-/)2W5SKW:UdZ??/X0=d,/N3IZ@_#9:B,07B](a0=
V/d^EeXX_.J:992b/RcN3fNSZAA@NL^FbaLd4Hd4fPSBN<I_RYST^)6:4-I[U+YS
9K/7HEPF)M=UXD3)FcJSBEQX53G;P-/()W;\H8=&a.I.&U;1UU/J?R9--U[=@N3f
=W&b8KD?cIPN=C:cf2F].BVGD&Q.-V:L(d&.IZ\fe7f<2^O7PAGO7d#^=43W27<W
\\_+GOP].>K?YgYP,8,0f)\F[#fJ@^3K9:G3Y+2K5U,TO=_0LMZg<_#8BH5,>g5F
EbG[RebK+CNd=ENaLT^J.08bHQGQNd&AM8MHRF\K(HN+S?3F&_@BGgWIP274e1RL
USGV1I4HeAVGW#BWRf,L::.8\?GGJdZ:9&cB_LUdV3;-GgU(7+e]X6(#1-?Yb-a+
J_d6(DIXBA51LGE40<09RN&P77f/B/9\J-aT37<c[.,bBTfO(6L:MW@;/896GBUL
AX9\=^75faUec/@^eYfJCBX5<I5e;1DH.-a4K_A&)34@AY43N[563II/_N#b_Q#G
E&)Ka6ZQKFC;<:>g_,82OEY:2g::ZEBH=I^CKR#M^M^,42AL>XH2aJ84-VK1H6R+
L22L6FF]7,#G=YLFO;L&49X0L]Tb-#9Vd6e/UN+KK0@^5:.@^IS9M?<R3I@\=e[-
Y4LcL>VW,WE4bSTe?^eU[RELYV7:;5MP>6<[dL8aP+SYIg<)3(+]_1L9CdR9fgX;
/EEKS[>]D<B2J7=d5BZ+Z7<>/NY->QX(03Z#UC(A(Y1Y6CS9(gH9O5.<+O:-GWg^
(?JMRG,,6BFg^Yc=0Mc-/+,WJ_5dS,,f.4][eG_R^YD&f+ET?D=OYHJGH#&cSeZ.
d+O_7E[>V\^39M[N>4+PK+;65H.f33:_Ade9Q3>CQ)JZ]]](^>E;>@Z[J\bE[X>;
U#NDRUJD]R[,C>XF\WM7)AAO0Lc\CN=519b4)gA1G]96H80:],dJO9fX6d,N0e#?
&WD4MVZQ,T(X90?(=Dd<4@<8\R)1<:7_agb[=C[?3K]2;OH-VEeWVWI/@a:93(:8
]WD1&BM?a::87UK\\J>TNaE9]H:F3(aEJcWV\]]5P>aXQ)KK@=.M,;E@@&Z2QA>Z
_4/^90F23C:KZd@QU^V:O+6Q5Z[(GCZ4,,6:/(0329NRd#e,:N0K,/R@^GR,\))X
-7L2?TJ&:0GUOG2dT/_3\.?VeU;C^N78<c-IfgT]XF+.a.HE36]5E@[5a:[NDD8E
Q@(6+>\KT(Mb48?>BVHegdC5^L)OdR0MZd^1:<HS8[FP<Qe.-R,UFd+&/e2-2FgO
:gc]?K2OK/@+<L4(g#KAfdNIKcOXT=6@bABeCZ^c[9M?-)PaHB,J3(Y(OAYWcEOY
\g#4bg:6aPc?#O1@9L2LHDacIWWRR\VCZQ<dA=M^L0fFW6b=9I,L555dOEdO+PG(
42R4VJRXSbTD:B,JJ-bO1;aX(3XU]O^QEf]=-9OQYM(QL9ZV.fZ>NT5N8Q^DUB[R
42@>_0MIM\>aCaAI_R&P3Z7?[6Q[<&K(?V\e-3#;2dTYG+1g6O@2K(J&d\0d]/PZ
G=J^?OMgE&(#NEQTZHDacGe&U?1662[V5ZMIC5daL_:2a<08V,H64@3]Q4Q8K&&b
AWQ)B<95H3SS&2aKDVSD,GXM;8=>ZdAI<<)NMMK[=]\;:#-d=&:1;0P(#K=<&dVB
-:Y?&IU_8+cB7(-E/b]E864)7?&7Q+K&;YW.6?28L^&OTJ;)6;cGb8S^GG.PE/gb
(SL]CJ3MJBLDY3gaGRe4J&_Wc]d9aRLYf9[eWDK_9gKHU^7E\EJ^g#HaXSOL-&\2
0g2I;MER5Zc5TZZ+06BT2KYY4db8&FHE+>QJfS@W#PMKAV&a+0[:/NDJ9#d^Wb]?
,:42>X([VY_]a;Pcd:U_<+4#HK,YUJSaGAY3/,]QJ6UE<#?=JP;a-B_]3E_JCE?A
05fOVH/A1cJfD^cbDc5&N9+586&-a6HXcB5869441G@L#)30E.Q]SBSU&DO[L<\6
.TE0e\6EXf,8Q1_.(/Q)@(@P^RK?Fb+YH<IFFLcD77XUf[W<WO_a2]fHYSBP_?P4
P0.U?@SF>b,Q#_KPM.S3IH<S2\(HMbWd>HKJNaTe44Tb2RIR>3L..S3F?_YScO#6
1^g8OUN.eZb24+baLJ/f:6P0^]4+4B3Pd&9b,/E,G;^4+0>-f>HbOY5(bVQD/UP;
MW_JHa@G#Z0a918Qf8@0<G>PK40K+,<VgRUDO>CT#6=M6^#RGJ,2NCH)=U-A;FH1
,<4b14:a5dIS_@>BKC;I)ae1WF[0L8=a(g>2U=K)<QG(Z///gcc88@K-;L3c]S]>
\&Fa&54RH-cQ7?J@2Z^VE=1XbeS&/PLb/EDIbWWga9+)=)dS+-a/3<<>QOg,N_-B
8YVE:GWYPW2X\>7DC)c(9e9K>M.=1:+PD5C44_L-KP6>.&XYJD-^X6?=6=][FcTY
aBO84\@/QPbWZ;eBC6.08[#4,=d@3DaZ>UABV0KT\NTEPI\)F&&[9bcdLeSLG/[R
4B3f[JbN4(447PBEVA]J?^#E\<aDa]CZB.PU\42;)O[HB\X_CM7DS,U;QX0Zd1>Q
,;;4L1W6eQI8@(]@I\1UH)3#..?VE>U<WdEND?X2\WU_?>f1;-YW[>a&C&1a;#ab
48gg][DgWUDOTc[EV;B3>KNQbgg-W>-\:7;[R]LC+=,0:bVg6YLW?RH<U77E_65_
?B2PB863>QI2JNAf].Z5T>e=WUT,5I+ST44bAY;b/:6[4S1:8KM:.L)dfY;9?57S
?E<F#L_4A#BB;S\FD_0R8HZd9dVP,+RQ..b(Y)TC],(1(aJG0NY/Wc6D)OHXV@[&
d&4-CAL(f/H:M_GL&TNCWN;UJ&P#:Z.?683NUf\ZR8D4&Qfa#UP;])->]XT2\)E8
HAPBH/C4Xa-.SN>EcY.-e[_e10/9&/[T@L\7caa^C4S4G;./;d:H\g#0M.LeK_AF
I>1=HOPH/(:]FJOEc7:S7B\&D38AD25K<WW0HS@BXS9ZU^aG_fLE:Ja)??([c^&W
6(IOe.E&L/A#6+]OB28_#Cd,=9W/CIaSW/5UYDEDWaNW6]39MQb+?>L4NEb]WDRL
Qd[W=+10cJ^4g_Tf<:YUXGV[K>@0AHa_CWLEB#PM3Y6B@+Yd^0?+?&NPf7/bEP/)
N9aSL>+\4F?e]AH:_G=IDV?TIXJ5R=L:.U_YbUZBaBT6Y]Q_<Z4/>dJfP^+<34Q>
TOIO^&gU/eR?[J2>3=fMRd#:7Vc8_fJ+.[WaL8ObdX<aAS=J;;#=A:[fHVe7OX/<
G>Ke40:bL<2?aaZ\O8[XaV4I?V?[P:/7-/-:NGX[a8YLM4]FL5ZX90(AR1^gd;T-
F17H)5:VcLBF9GMV#SbC(46;GGQ4=YNDILCG]N^;b0]Qc&?LS[[Qbb\<aLK>YD1[
^G@@3Xb>MQZ(Z9&F<5WR?L6He\>=[<^(/JfD2LcE22>AEdT&U(\d,f7Zd5WT9_cE
#.9Pg/RW-X=)4.[(Vca[d;[;L=b1HW4@GTO;)#-+K5eg<E.F>&S,W:c78^B]X:2W
OEF/?8OB(94;CS&L_cGLJ6B/E.5cdfcY;cE7+/I1-:1b0E&)+Bf@[R3d@[efHM].
Xe8PL[N581#0@E)R?<,OL8fYKa+4W1baae4P/f\15T3_fE+??WY2@d&NP7C\(JD\
FH->??5U.SG&ef=0.2>.=Z1Q?:665\LLDgHKc.AOB-DV#<DK@?T(f<J1]5;7e]&3
Pd4\2PE4#U54a3M,^B>)\-^C#_FC1R5<gSA]N@X4bX12<QZ+KGKN[cI3f475g.K6
N,<EC2bQYNS+\=d3015C.SXQCOeW0e6ETTP8a-d9/P4E55>9H<JQcGAgQ<G(\ecK
\X^39]1]0.M\64SC/TM6VCU/<S4L-?-IZR8]e4,0#=AQf.JE:Z<55;;d,)2-F98=
-5DU3U_<RaGfF0PSe(GO6;XX4]dd(7TQ&V\JZE\X72(7SKQ/7J=MO]LU53SOf&W/
J(T/D1)d>KW,&(6I3GI>cS3bRJ_5(47.)92IJ=\\JdC)I07a0::JI>Yc.a=g1<-g
HAI3RR;,Bf;2T<R9/],g?G444R8X#<aR;\\5f51CKNH^8O01MI1E.]=4?OL]2U@]
dM]IZD5DICZ?J/AeLWTg&>H7@JFeBJ+a#QfMPa340@Uf0SbY_f4Hef2;^T-8U0=G
b6(1=E//g7=6T&JH48;76ffVG^G]0L,)b&F50GXVBB_:Zf_Y-fdd#R@P_O3Ya6)R
BZFBSB:e0&N9]8&GIQAR]L1;2SD=98X4F]2ga<&OIUS@/HKf[84?6ZII1D0[2cKQ
eLQ?,dQ)c-Jc;@\beLfeN-XHI]16(\A_&:#^[)E[gGY)C@B86619318WQ1e79FRH
CHV\f^L(XdbWa]C<:#JZ-0F6YD)@]M?5O6OCZQ@dZ39(I(?/MQZQ6UBF?gC:KOC<
cdc@9V(H\-X2M3GLdH\U[]?.3A)cFJSO4PVQ/J@Tc^f&^?EPT_GT=GK?-W=^4&W@
1+64Y06^V45#SV1<LI)NUb&EO-)Y[6FTa_ICQ]-+P,#]7^F6@dK3N7OVeQf39Rd^
-.+SSYR.BP.6]Q/7)=IaGVJ0[+&LV,O-NN]gBKY[d,-\^Q)H0G8O:WT#gZH/d:FK
@W5M1b;;)_JN((^SDY6P>cRWA&K=[#F]F-,5^F5gdL4([VbWU:R37K7RDCK]Ve_8
aSI^e8:(1eK+51QKH3(RV0]?9/[<&K)1d@RR7HG([(G0d_PU</2C+:0CKJGG5F53
b<8+JR0MfI0&ZC)YQ<KK?]fN8VCOC[>[V=1ZSa,K5#Aa1#35He#]QK\(5AS0?#8c
;P:SE-(#\JOCLb_/J<PI)<+9\0<bTJ;O2ME+W[D1BG,&Z]PVTd]40,CU@R+S=G4B
I\RN7HR/NOVaeK;EcP,PKcKeLU]K>3@].S:P?H:6-e^g3^^V_-BdNW2Y.BXFBaG[
G[cIUb^/,VVFb1aU_.d\OcY+HU_K>eRU.3Of<-(NNQ3_HY9=;f=QBS=T0/7=&&@\
_C5P.]0Y?4Lb6=N,OF([>(?<7B_fc2]<,;e54ZS:@UX[)/^0>J(VSEB>ZQ:K,8Y/
\>RZ4N3O<?3&Y^2S8ce8JBFCfF1I.9/GGAaM/3NSBF&8VR,S=-(<TX\=KJ(]7&UC
Eg[OT3@>ODa3ZIW)((E<02PdMcPD;Zde97M,K@?K:OCS5Q3K7S\OgdI7Z^3c42]Z
3fbWO#.daS]eREJXLF[dP,G3D<#1BWPgf.3bGc7KP@Q^;XE/5_;]4:fE/dI]@^5f
,c^]d:-(cF_/c#\KGXa)Md@0AR:6L+J6-45RVL4UYUecU40?0Q.TDU)F1VZbP8;d
Sc-R_a+LYK;\,@aQbL9;TCGZR?1a-?:H>f(#C8I@b6:bfVCO4ESCDd#:_/<5S_Tb
(Y>Z=cFaJ^W;@4P:9[=1@&;8_L8Veg]?LET4]OZKX/FbKgUK&?,Fe(d>fS-(Hg[M
&GTd9OeUS>5BUeB(POGd(0U?d4eDK]TPV<:bbQ(44.^0X=PMU>0\EX4?B5aBRI3X
]HN/@=:RJ]c1L0EWebcEZb=S20(E^F4.#fff4WL-#.dI@QE8ff[<8M:2NCTBd6-.
?;dfQ6(:L<f[7<?6?KUPAGB.IK&_WEQ01dQg)EM#bW++4E1Z+>7N0eMRB:<U\X=?
D[714XRL9<(KcKY#L#[NM+,-\>We?Z,C/HV]SD[Ob5(_N#E0Z3N2,:>B<4\-,0[,
<g[[#dD4DeEb]1W#8ZDReU^4WP2L9ZU0WPgcMYI;cMBcGVa:]&[W:+N<AGU;J5a\
Gc<@MK,bLVZ5=7[(Fd1CW<BOb68)JY3VaNQR8bfSO?0f-4VC2XED;)R(J;.PXA@Z
W;LZA0fa[E1M)LP8=:]&?9Y;/#[d-]#MFZB6Ic80cC\:>ZN<d=<;KO6[?HXIK@\1
bP)G><(ZZYKPHF(QA2PHHX;KB;]eeV93OG?Id+_ZCGV&3I\>ON#+P?S65(\-@]8:
-7[BJP00KLZ(Y6DM5&BKN9O+JG[F,F]-:eR7M107[[1Qg4KS:?9)-0=4F/fH,UXS
4TGf>F;IPA/[1WQU_:F^FD(^-VfQ0G#WP>#b9O=8e@O@CIF\JgbAR7c>+e^[2.N>
)@]DY9N[Gb7ZN0,4ITd?6_\6L?Yd#ed;^@LR6Y21O\(7PJ7X;B0M:MT\DR#\cJTS
VEW&]B,[.Z2b_-<O?d1G9;gZQPRb=TQ]2QZBY>HTHD,S5&@He.@>-_VC7R2FYL3G
gF...>U]6)3/+O,gaGN@#aQBCgbS+DfH1dG7&UK+A)]QC6=5-B<4c:<ADYg?F,a1
@aM_:Z/@([gR)I_RL1f2U<]H+EI[IG&V4^TLC/L6[42..d8#T6(/FgP\Z.b:#Q2U
AG60>LSHN-S8[U.QUNA4eegVbAITK7FGBB6DNdR5P:7,N1XLRcO4We3LY45/YN+@
820;6Z]:\#)3N+K,Z7d3bKf)]_FMRO]&M.TZ9K^TGV8,JgM-BPY-_UZ@ZH.@gM8_
-XIa8PC&0HaZ<(SGLL6\FeV:ZP+NR8[D<6FQDAE+CN,e+=SK8WH?A#LbZ4W:9=<4
HXB(5ZHJbC6Jd3-8A@F:@C3cC=;+LE[(H;?Sa+A;1P,\W?BL,XN2H>F]I9OL1PbI
YSY?=gfO7?=Q#9cg8Zg@QKC;;IIE;W3P(Ca]MP.bc5GMU,Q<FLGaOD,,I3.6Q#^K
fG3,H3=?(]/L(<YK5462:FT#8b,3^K0ANDD64DY?#H42IVA6)^gO)Y@gCP_)2FK2
f<],H;3(BHECc-X,)?ScN/LeFJG(5X4gb\UPM[W9gNg(SO#EAJb;QX:G^B&FK&/[
0:A>QV153)1&5HJK+32^U7#K-PE6e)M.<$
`endprotected
endmodule
`ifdef RTL

	`define CYCLE_TIME_clk1 4.1

	`define CYCLE_TIME_clk2 10.1

`endif

`ifdef Period_1

	`define CYCLE_TIME_clk1 4.1

	`define CYCLE_TIME_clk2 10.1

`endif

`ifdef Period_2

	`define CYCLE_TIME_clk1 7.1

	`define CYCLE_TIME_clk2 10.1

`endif

`ifdef Period_3

	`define CYCLE_TIME_clk1 17.1

	`define CYCLE_TIME_clk2 10.1

`endif

`ifdef Period_4

	`define CYCLE_TIME_clk1 47.1

	`define CYCLE_TIME_clk2 10.1

`endif

`ifdef GATE

	`define CYCLE_TIME_clk1 47.1

	`define CYCLE_TIME_clk2 10.1

`endif



module PATTERN
`protected
?N\;Pg:F[/7QRCGWC)\^b&;^D9?-61@YO>X;dJ?EKQ/)+0,>QYKO5)\=H5]14,_C
CQ]UDOOXJG)+(:1VCIVeFC,SD(G)UMMbND<6V,\O>,0_([]_F9=^2d2N)#0O>XH<
HCV0)5:QBQ&NM-)]^@I;SX+IC:bS+.F;==F&ZH3HO3];SS4F2\.f[;G#,c/,eWP&
4=^/^Z:a?5ObGS5D1OP\\D/>4M&=d6M_)c_/SCJ,4dcWGMc4T<C9DdK9M@PEJCBV
[QRF^YG1[-6ReZa+9HEaX>QDc^#AYg#9H(PJ(/9\R5<8)@Ha>[<F@JZTBGG_7@@5
N6>&bH87J0OR50Je.g6+BB)=?0?\TdXEC&MF4CU4bO(43fG<]IZ5\=MacYHF&F#/
6TSD#9_\NgE(W6L,D-MaIZ(R5AR4GX^Mc<N26WFS8ZMDY-/\6IDaXR&PKQTN5MKC
&Q?CLFP0V_68C<.Q_C^IO1V@6:E)\C^ZYXHOVFERH/>+-CZ#FfEC8bQR/PTK>/Ke
#OXScZ=dB<CcN^G=4_-e@MEAYL(gLX_R3d,2AaFDZ:.0)9Ica2OF.</74)C?,.@\
X8X)4S&BIWZ&Vd><-ZQcFD-;<^GJQb14<,).K>D)#SDI-4?T\P(-=2g;(_OH[H(g
f(KdE<?E<=\d_<a.FL+\PG&MOf7)3SKNTgCeWO#;;=NVL/gZe4gJ2-Z(FM)LH1SW
M/:e[,f6eHA]T1L#d&V-d(dJS@W07U[\81=ZdaE_L)=9F3L&,N3-#E,K#+6P3SX2
4X7a9GE/\Y\8IB?g?OFEW&fD,^/@TZ&.+-b,T66Mb\,/T+BP0^PPQ&aSZaf2.]5X
4_2R>F-aG-VOS9D7EY>F/fI_:DT_&PK?_1S_<CQ:98;6RED^;FD@XWJKAU6@EB=2
Ag+69-T\X>?76I?ML5>?KG2H1]BY,>#3E](HFA6NQUE/64JaBcJ7@MZNC(8.ZZX8
fTC[VBV:CG9fXb71]QKN;<X.-a.>I)ED:#JgILYFSL+A;@K[T?e6?SXbGYVG3/P&
<E.gdQgbPW;17Z3&/X,LD>+BgJ.?[3^./<J8KB2@ZVYd>AX[T)Q&NZLc>60WMBVU
+5HJe8VZGQ4Na=Z.&/&Dd174MGge+K5RC1QH[@CJdd5]YZC<K2)9T7K/Jb)=TeK=
HYM7^2[PJV_3fTQ_97\096-(GcPST^4R@d03;9Fa?_0<GKE&092S^dS@(SBd=OA5
,>.4J>U;e-KbH74&YVe>:18Z?a40-KLUCH[_ECGRSP53g1e1MS?G(L)[<8fVAIT1
^0@&:M>J#9d5]A7N>T+EFLDb-&D(;gDSI?ERX_9]e&V/U;N,]K>EaLA7RT^?<459
G,JS9@:JHc]?[-?AIDZK:-1bAa&G.]EYcSW)2,Q_IGUU.]Od9VOcf.O1=,bF#acY
J5))V2#7b71GL]2,V[KN9.CYcA@dI=#1D:<6HgY)9^:7A)Da4a,JfO<<MYIF[:9V
e1=(ODU.R[)BWD7E5DZB02W#^LAN(ILX>WG,[WId>OM?;-XJZ:^<5SGRb\LWI4O7
M5CQ^TO;<Y,0TgG.WM0^G_PLJR,1FbT5H,S9YTHT]=SDB[9AY;eJZ2TP<>G[W+QU
G,E.Me<>eJ8K[eZI26Cc5cX:.4)1bBHH]OKY,UWIDfLV)fg@Fe7V/8H-2-E9JN7D
B/0?,V0e&91##9aRdJ(HAU_,#Hcc,&_YA4&)48@O]9??.5IG5^Pb)14b.&gK>)[f
.0Xf-:W+4agG^@^cKTKYBCZBZP_1/gg21R-Jg)S1a#e7(#5_,_WE7eg(cJUI[3aM
OI2U[W(FR-?4\9gCXI(1d?d]S[bWY]c/J8=Ca>54Q_TdH>8=YN(=/MKGX(NOZIQS
c4?7QSZM-=)O=Y4AJS\4eUUF9;&+<6&Lbf+d\AK.UF<QRQ[XU73b57RN80=,be_W
(H_P1K8[6aCDa1)9UCd1cTZ0)^ZNX051(XKfb?(Ic5)BYD+NTd4(_)A=HYLIZWXd
,&PbRF1g.=G2bL3bZ?OGN,N0g4-457U5@O-M(MQNUQ7WS/,?A#OUG711,3dJ)1PY
[dA5E&/e#C73X[.D#Q29,[.f6#G2>MEZ=Y]bg7FdJbNPe>bX1FSWTCG>+MJ(QFY)
VT)O]\LFEM7_af^BD=RGe=D:41S[_M25eQa3fbM3T[6F@O8/YSAgTNI#deI[(\,V
[:/\-2NgNO-.T[<<C4D<@H830&#E79S[3^E,d3QeR7Jc8+NK>d4M:\1)4BI/:4<>
<M\)DZPG@W3VKQ:&JBe:W/D@MD5Z]Qe4fa#\WGI6fEC\S7=HC8PU]X0B0O<]6).D
6_:^+7c+ff9ZfC24>8OWJ(;Y^NgTED.4^g0<Wa?TI.d5O-JS)FLALEVV252R&_77
:]RZ#6OI14DIX?26E0dBa40HHI=3RG0d#ODYdD3>+9:U7BO^#b(cSb0=Ha[9BXZZ
)8f5FTGPeAHcZ=U\WSAf8I>J?KDGLT\:-(dZKD)UC?I7BAc@595fLG?IUQ>IEW=I
@]D<^B=+DU[d[MFY\JUDe&DG.Q35PZY<42If,NBO1dcF=4=234,(R9H=1R?HWbEV
)O3&29bQ-gSFYFJYTYFNL1Ue<GPIV,]0DE[_PQKZeC@#:)c\B/V([#W29@-P:::,
eEK;g@#VID^/Ta(SNQ-]:,?6HcF)?9I3>A(H7:eC9LI><I;LY#c))?B^:181OCI9
^3ZD>QBU,FBYASU&B2/)>8aFbgL6//1_>A:Le1]EM]F#.7O\(YT(C7Qa3T&YYeE6
S1=+\I3?^a_C9,RaF-V<D@ee9FG^38C/]1Y#MI-6OWZ6aH]Wc:<-24F?W06)^A2b
V)deD7O,1B;==>]:aBaG64::]6SK+>-/ZB1N9dX>\S[4CL.WRM7A9=K/cgNMX7JX
.R5R(,Y]FHdcg.H1bQ\2H?ED;J7aQV;ZCA6WQ;1XXV-af#N<Y8:e<GLHL<]KaIdU
Z/5VW^7:I8+UI>2e/7K@gg<2&\6Z4;e[O5,/)^))8?<GP.X4BS+:+ad[g[;O\L>3
D7:M)Q9OfH-fg1cV#dB8YQb>+[fU@V_EIW8^8E-P,U)_:2^?aF95TXb-AC(>L#aX
SafHNVcF_?[]NQ^fRUM1@Kc6/[:c=UO&)_Wf_cSQcbEK<S_bSW&Q0dOX<da?B?;X
&c-3T<BW:_@W(/X4_0/3-D<S4NC;=1O3WF@^McNKV[6<K304]URf)JMSc@/)eQ,7
-5<><U9Ge:S8<&K(6a0)/8_#6)Q-<geX76EPNHASYHWR.6K)^dJC+NQO2JO8K]1+
VZF#0Y#gFZb3e6+4Q;\30b\?@L;(?9F_d+Y0B.f29]b(:N816aRbUDOR&=:?,8QE
?W+f6]YI0FNXJ5(9.(WQV&KM29H/[aEA\8b0:S[-G/R4HS9+0576+L\TFaR3?_Qg
>@E;M@-XT=MaAZ\K8LW0@e759EeX_478)D^_17OfF70;+Y=].,3G55]f^fOU5I\,
OH_d_B;cFNB41SI[<SZL<&C:Y#E^F3[;O1D7;D_)g[X=]SS]>XQE=O4GCJ4dLF7#
a>I:MT7N#QRNK[A_I)&^Sc<4G@<+),<W&WX\E8[23N#1Z<S]>1ZHd+4?D77bOTF?
_d(<7_5J=T7f-d0,G&M8/_]7];==C\@]J^D9_[R;cId#>I(P(&W[M#@_NA6/HEg@
M(&cN2QM^feQF&2&BU:cP=3I+K9[+N)7Be5(8WMHbR;M&a]W/?W0d<I&UZ#aAP#U
0YcY52JV=)L00)>QXdLS#&D\e[\.B7;S=#dV&9=5RaOG^Q0aWVOV[bV@QNO4f?ZL
^&LO?.<VJ#X1L]HaUZeVa>RNTFKc)FOFKW:SeF4-NVA<g<QUC@(VeS[bVO&S<QMe
=D8M:aYg4aEV]_H,X9ONN3D>e7>MVBD-\ED62N/GRD=UB4@FM_YMJ3[[KWB2RYJU
A?;C;CgKc+:+TSXM7P]8#E-1SGXMWFF-.7>LOfMG2eI.T#\;(Z=NVc\+,JD/<:[\
PGCHJ<&/01@)S4+.I?_=0LK+TP#^9Eb,-:@f<CNaA]@Le,\g>B>8HEXaeFfMNPeW
ea<a>Y_?4KPRLU6K3\^@P-g^N++Y=1Hfc-Y@Dd&^CLRXDdS,NU?SI\VBe-AV_0I<
O8@BQ0^UQ1=:>g;eZT_Z735ZRPTPH\FQ,4IN,7\_]>)Q9bDRa?WYD5].:=&F7aUd
?0KQ@O[Q@dRQFMLc7]fg/,ZPLc,2J-(6eNBQ&g7^ggcL\dPG[+E@I&V5Db8/]3:H
Z_#?#<^\]B6ZHKU6L5)@CCFW&H2=2(YT[=UJ,<W;bA54F&HNSQ9).a:[^/dL,1Pb
g]UX>I>V[A@6/_?-17cKR<RV[^@fQB]I<cJ[W@f8PNgPEQ9R12@B;A-H+Y=@RV(S
6cX4fG.^.>1:^T\5G1gN_A^4W0dJ5-eLTQJ?b;MWCALL>TYAXLK3_P#5b3B^Ga_T
Mf<&>F=&<f?gdK=)GW=H_IB;4aD)]18F6(]Q+#GX9IGL?.3cD2e-[+Q6RP57?Q,#
@TG@f&acYA#JB6?_#:SQ>,/fW]]X;JBf-ZdP46f@7D91BK3LM?3JI.SWV^1Ag:6)
,dY>7gT/+X<2bOeL8K+Z9&Q^]ZPR@08TaR94XRQcUgG-SMEVT[,K+#9(7#\a?+HK
\dNaTS/C^J9@CLH&TSYg/#\5B#C[0),4JWF08YAbB;83-@fWPDa5e;UfE5&I:.Y@
T6/Fb8I13<)c_[=d)X?Kg@RAE<f[b_FeQ3J#[faI&5OaS:?V/=(-#(a+[:1=<;&,
S)CeK54VA[Gf9[I3XMPF0c#Q-D-D-9F#:[+0Ud=21HaBR:A8Z4]./?5J]JG,Zb#G
c2FG-Bc_&O<U>NVCX=Ga\>FUW^,GC]bBBb_;GHU(MAPJ#K70beV4Y[>]B_,[AQW=
/@3afO,,U^L<#MXQB,b&?F/W90XF[P[J2=gTLHVOQgKT/PNV>e93-g5BbO=JUX1A
(bDUbUOFP4I7B0W-I)QDf]-B/SU(Q:/1gcV_+]?6VW>adNec[)XY7C99bb\D_?=?
V44eJNC):A-R4(ECXA79-KN,7)]UC56^6<=.WB3_H7fL\g64?2[EQK+#&)T]HaI;
f^R@;<5AgGYDW,B3Z@?Q17]:G[#PdG^eC1X&?6dTZX0WM^Z#<#7RfG8.CVdd3;_N
5?OK//+2FT@+\Y1dGTD-/)(;8=<3eQb#;EYD15-CVLV#5(-:F8Z)-TO.0JFLM8f2
OW732B)CP1I9?8d&-2-Y]TFd2EBF?R[GQP;OC^B]G78,]-#<T(W6d/+f@5741C=M
Ug-2Y&@ZgGJC?c38aY&\;\G6\I:KGZL]V?[d]Z_=]XM158L(Ze+T[&:YO(V.JdZ.
H1E4EM?\bU7.dSReF/NU/CaMXRX6.I2M=>K.-a\0,O\CU7/FG;JN()::7<5\J+,+
:XXU<Cf093:_+;KCH>Fc>C4D5Fe5Ba-\(=>=5:/7WVYRP#aTReYF_Eg[F+3dMe4+
I-9Je)7#9c20?2LZ>5.K23Se_b_a#1L+5N[9,SWO)951d=D,04S)f=B(d@B\H#K4
M<MfAgWQN0Z^;Fg(BW&.1KA_dG-bcI+K)ZaI:Ge[0<2.CIK?7CX1fb\eGF:QY.^b
VeFaG1UFXE,H^Lb(.#GPW=ULe;5_<XQ/93aK7gcG>-1agUbHR9-[U>LE\LDB3_:X
?:>dV;^>+3\a99=5QI91WSb\6PK)IJ?Z)J&>>:?KPQK>b)2Cg;=:W_9ESM[]T)?J
W7.bFYQOb@@AXd&3D#-,&&d[UO(>++Bb2YGFN_/)<cc<9(c@b,18A@:aV(fRb>;5
0?\XIDA[^0&C;VC#\LK5+Y8cO7B,2A:W;1bX>,APREIWSVUBeA?.Y?f>:JcgLA6A
GQOY5(D,MB4a8OTJ?_3C8&>9^,K9OcTUGaCBb#OF&^9QK[NJ&9Uc4,(?[,RX#83c
J:Ta2B9DG@=_#G^Y3J-XZO;>DFS0e@8J1E118W=^H;ZB[+b7Gg(W:1SOBW,f@ZgR
C+CA=EN4#Ad?37\OMe>,M93H221N9G4,88(+AH#;PNa<dAG5V-BWXISfL/&]ATVI
df2:]1WD783;c-_gHRHA?7aB_0+=SQ^,#O2fdF4J[W+QFG6Y=]09#c]e/=@QEdH@
e<0P5,DHF=D,]@NY6]2,@QMc<+,<3.T69gX4>J(31?5^gI2P^89)N,]ZQUbR?b-f
:WO7=G6<U]1#KQVYE58LLR_-ee>4VQgLTH[cZ;>CN5+a@[1Q@3_5fW0/(bf_DYT&
b+d9RW=;.X0>2#YXN^<XOM=a)9_KK2[M^QTM?f+&dd@ZcNI,KZOaW.D/.d6NBPP5
gBHVQ(A_76-@=GGEVE#D7;P1K?454d+NbT05G[dD8&A5fY1bWd7O,8S#.BC8MPe(
c;,WI=)(IC?4,4DSgNA+[;=F?\X;TC6^J^Qg=5aOdg<S(^6POV<Y6A0+J^D&#8BX
5QFWOY;.T<F/+_AE5]7EUg#^RRW0+e1+0/E(49M2c+A=F//]<AF9TY=DWA<2T0#J
IdOcHf@#?:PUdIUd)SWL+H2C?gZaK]A0__[#ENcb7K>/L?.]D1e@5<f;9-05CD+Z
EW(eKbKT+V#2CF,eVN3J[B6R(RI&6YIOD12M,[g<U[Gfeg5-?d/I/+BUMJd\gGJc
:3H&GP^bKdWE(_+I75X)8,2BICK,GJ?_)0<=D3[E:9J2W/J\^PSaScRM>;_+(fJ:
eEU=(6g)X@aRc#aH3UI(WS[Y)f/HE@@_cA3a>UTHL\FaZA2HZ1-:1+-6HVY4(f3A
3PFF&[AXDVVS=E+F&@2fZ#==(\:I(dXIUY/JeV64_C9QA9I#;8+dN-&BS#Tg58N3
HVNED.O_E+L,5VFM?I5#C):T<4=UK)(VLD=J8T88QDCP4[GfW3TSG3US?;&V+H/+
3c_)#F3HMbaYD[>LRaH[#KZ0VJ[G0^)8dK-ZW[ff5PbE:5U;g&C15<@aDcaI&cAE
1QSTHG6ERedB>A1)&?:JJXcH7eT?5WB>8KSO]/9UYG<REOdb6?8Pb:0..&Sa<Z5I
BQ0O,3GVDOEHDO5c^JK@_SLgQ<<-E[3,9\3X9>aSE[IDXBc2O3C[T(F/>N6aR5^N
6BR(AP6e+7N3D6CA>V8<a,^#Y@U>]@2(^cG#G>0<9d?A=1YYN@O98@J7+6fb4gMG
AZ+XCQ(@_\(\KEN5^fAK=->Ib.C;/WT8\7f)IgIR7-W/46SBN9-ZfC01GTcV\_Z:
;G)Q@W.:F3ecN?+RBVXITE?REBY9Df9?T80:TUHZ+_\K6(HI<S7Vc/Wg(?&W:-Pd
b07Pd^.(.RU\9D=OY75:UZ6fV+T9QL]aLOe8Z0D(-96#VG:^#O0DEcL6>J?B1)O_
g:ZfX]b0)aK(#]\S-WJ@]Ig):McFJ3+eHD=48R\2.X(aD8NJ;1\C38?6A6M+:F/]
KGM109E#3^g?Z[\ZM.TE6/,a71:@-7Oe4^Q5M#I4I]R/B0GJ77..4M4d/_),HOTA
e3[>DJRZM,/Q[<IGQY0RJTbE:>].5QfN7A7&BV<a:[7;,c_NVM2M9LJBg@V<E^P4
6-&--1gbA3IJFgS]:]RAb9GO@S5,GYFIJaHaIIW)ADMJW)D1DbQ1508DbdLMH[8E
TV:VH8=PLL4b_+BbB4baM;fbNMFX_@VV9:D6W@RF11faE9Te>&Ud?eBfI,aVU-G>
ZSEaT6/6XZ2><LQ#a=V5V8>,=c1G7FWUO:A+7>F39<NBd)HR\Y4Y&Bb-1Xf)Q>g;
A#VQVEQQ0bXVZ4I-B7MZWRBJC;b0A4M=b0\FecZ8MS&:d.L<NLf/)T/B=8/XOd+f
WR9M#^>BVAZ_UJ/F<\f=@ZQ.0;>2[,G@)(O:X1ceD.)1:]FL8@PNJd_P[/-dJTEL
@&YV9.be8^U?HTWb7I\\F]N>,9UUFFf<S&-Z1-CELXKD2@8dD^6/XA1H@R25>][9
GV8d,QI?C&fA\c),X3Wf\IHJ_+B7,_.:,5IDb70)Ta)_)JE[>;T=_^+BJCA_\X9L
XC)-.#W1+3,CRg;PeD:gbOT\P\E[_e@>\a_._Y28UcG:Cc+(/]Q8LPV[:NMETODZ
W,a,--\7=9=YC(_6O_T[<<(X.Y\V9G(=WaR.R<ZBA^^0116D\gJ;,WH+RfG5&J[=
G7Kb(46]^fG;E8R>G^/B;:,29d)Ze8AKHK7#:Cc#g_6+>;3?VBPcbEH(XGKf)PdB
X&BUPI2+7fGO_B,:?NUI#RSFK8S6/^3E+8IP05Lb19N3SbTdN.H)cJ5P+HYR5G+,
a6_IFC<<AWCI#eY:Q<XHJ]@RN8<Ya;8BcbFI/HHCHee>O+:.e4J<R=Y9Rb3YV(W<
V(X[&cX#_YJ](,<cRGCgW&S#f\fIKBe^+\^g+?d;2R5]YXIWa@eKa&)>M7.Q#FGE
NF.]8?J<I;24?(GOAEAMC?8P\IT+)83e<=LN)E(EY+f0[7g90YV5J3J<gc[9((5H
?a,>g2&#;6e]G#dVN(+CJ:[aW9YCJcU0P3d^RPD<>\<5O]7^)@,7T[8D:Q(?5\L?
:KbI;S<71-OU5=BXRH&?9G6aDKTf2G//1gF.>8#-:&Q8ON605Q=]9VScB^cJ#G,@
)a^#V833A]6GVE6,2-X.eXcKEL=#JfI=?9_\f6FL8M#G70,CABA.0TOJ\]<d8=6)
KL.5^S2>KWGA=\A-T\OO_(29)+ea@-N_EG0S&b-1TG_cF:-NA5B21;#KJH+&e0^L
(fSc_BMQ(J3SQ.@/(MJcfWS+\f(91AXOB5^C#;2/KY1=5ZId66SPIG4V_?F.(-CS
RI.62\ENJCNI9^#QZ^VS[(+8Fc3Xd[JIB^8_Y_0\:a+S9Q)Z9@>&I=cg<QS1EOa]
&#Af.HA[#9(A<??A@2[Pd7.Z)G\\_fV[V^S6Ee&C/21D3X2Z]a2><,PYBOB+EVOE
?>.TEML<LPBaZ)_B<7;XI]ID8\8_.QS,5LbHU33=6Ed<I&1AK>UUP.>Y4Y9/&T,S
\+.^FS&B3(bG)=(XaDG:]3.L/bC)0C,W#OgKV^dPNDXYW>PR<]f/7Z6-,<DM&\--
3M-1^gg,5(:+GV7^gOA6Oc.[U&):9A.eBH@5N?6QD+3??<P?TXF6.CfP0HLa_cDK
R>@Wb>SeO+QDPX\d(BK#f1[7(aG(OV[Ldb.R^.\_9)\D7</Ib6:@ST^Xb&WJb-B\
G=&@Na/7U-5P]9_E<9=.fgb-1Gd=\;OM@8^]&3B1+.8G8IHcbYa=eee=5^+PQP/>
N]ZN&(C[=P&:X\GZ_U[SSC#<HZLYObNA0IS6IN+JPQ_K/;MB>>g?7?BM(;dN\^2C
WV4#RUO17=@;PD:R?N43X?YBX>K)OHHaG\T6/#BVb.Ha+KZ:C)S2Ra)GC@d\7=g(
^,26De?GD(&T04f=2.RXZT.Dg0aP)\g.8dHdQ0H,C_/-\8]dZ/cIX&6<2e\cBbe+
V8EAf:7b=I2U6IYMdX-YSS&^\b#UX>^ObZS0HeWA[;Z6UUJ3#(FDH#]>E5eV.L_g
g(M>R+1FPID,b+D^3\C>WSZ]Sa-[=M._&GB1\;LI)EaV.-P+9e6T(0dUA18]+FB(
^)TWcK&/<V98La.:?-&Za[]7+M/fPS[b8;JAc\6W)9<Ed]8+);DNH#/AA3;O+[TU
bSTea]d(9S5=?47dTK(2ZV2[X\0Ib5F,R5bM]^:Q0bdTLK98RNNU+W(@Q-^,<-&c
J7G>L2ZQ5A8CaFI,)W_XV(eD]B2#=FF,CS[Y^Fa\5Hf?EM]G2Y-UN&I&_NG8KO-1
_T@_\UD>B:DF2C?g.@X]YJd1gP4>KLV60#V^<:Xf-\4DfMa@O9H[&/=b,N@1_aO0
XIL-8]?&]6BU.]A@C1(gUX1?,^-:3.>]E]a\dB/124M0+E2.48?IR>dT2^7-fbC\
=2dKGEMV\bW[abEE2M(1@@W-Pa@UF[QP5>5(HSfU=.XZ:cN-#\bIF6:a?b]J)^9.
3GM#+V:FN7VD7<)MQ/7\&eR=?8&D)B[@K<;U;[Y?2R6PPMII#7[(d4V?R?c;<aFZ
0-0F7H=DS#177:+&PRg>X4>?41@WdK)7MPV5AgRS:<6.0[F?dNM3Q^<M9L35(OdX
?:H8a&/@R9_W+,]QK?:W/#Sd=&WRaXK<;=F;N.eCa]dKMS-d&bB)RcVLVg0HK]6V
IZK:G.^9Deb6XE2Y;Q6#20YA\-<-SHTF]Og(d#>J&K>GM32QXcDgO-X[CdP;W.[F
NE6>I#359VS=^(^c=NLVNI?K;<5/LE:ZMQDe;<;\fWAc3=JKSaE@R)2WO7<DI]=P
e<0XE9Lef>U2B_?RTBc[4\:AM_O=/7]9TVRcYA<cI>KZWP9/(A_IaS:aVK/<R6(I
D91^3RO-S_C+M27bP.B])a7\=&FG8D@^-XV=H[0dQdM[<IRA/a0(>/1RX3F?V7VX
SN7deL@bE9N3L70D,Z(JcJD8aM2f@P\XH3M3^ac:88:1X[HYKdbA&ec@IK>T)DDe
\\c#3dAVFP<9c.^I^;V8c_ge20@ZfSJOg)A35&F,YfV/a?.dGb6YF12KBLAeBUQa
DSG]3&Q:UeCZ?ad\<SN2JFURGgR?,UZ0:LJ>]G-##HNUfORW0>[E+TC8@;CC<0.S
[a_J,\)U+3Pbf;KdT)G@SO<+ZIHIZbQ5<_Tf-GZ_^[18[[/(WUN_V,OEET+C(BLD
1J=f=bO7@J1eg<5-_TLES).U<d@<<]E#V+1(2N>Tc[&2+:SdQgK-/.YKU[cKR-7;
^=6La[Z[]_F6[PO/Q&/Y,EWL=1]S(Q9E6FU8-XW>E&JHUO,Nb&2OTcC;S?HT6gJL
F[F6_58T#6\1<ZDFN\SBS@M2C7JB7fU/-g_B38ZF^SgXT8:FST?Re5:gL5UXAK2O
H1FdSD/+R99d,.?I:gWQ(L)1fR/#>7O+E;NH+9=;J[R-B2#33K^ZZQR8+g,^H+[M
Ja2QTWN8Bba&D7=e2/J:)0c:1LDU?5_aA@V76Y\W)T_P3K<S=3A3<C&0Z#HZOI5>
:T&gbK(cB=N#ZJ;.=gI;F0c_8Ja>:e90/A)6L4BDM6XX]SgVc5JUbDI3>?Q5/Q6:
Ka>O@^INX.+ZE=PG1OX9(@OONG8M(Z73<??F#B=7)K.d?FPc7V>)FX#L[b49EW07
8#faPe,MX<[f806Y79_.NTSV,Y4S/2N1FQDR>46ca)aQ2^^d?]#[f=6YRO42_W]@
[dEd,2-M8bb1S]\(e&Y9c\5dX4I&4Eb@5^U1V]T;ZR^D93ZL]^[)&fDK5VD?.2S\
TR.P<Q8\e;-1+YP3c9fDfe(P=KA]LT0F5W)4WWM5g;C1=/[N.e#,0M:0-(]FE@72
:H/K8;A_(3IJ.N\a6ZC?PJ[R>6V]7c0fXZN-,DHUQ7>/2.9C)LY>Ke]@JV,TQK/\Q$
`endprotected
endmodule


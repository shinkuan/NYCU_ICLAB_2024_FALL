//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
HQe7vrNcLhGScN2rFuOphYXIAZXlJiWDRA+6CSkNzNVrDdv3wCIjpNEf0cWdcRON
EJpTJFxeFxrlFjguMMWrpfINkEBVv9SXatmwA3lGGMsOWe4kCv2K/frZNOTgE4Hz
jfxikra3BVBL4YzL3TrWHR0Ta4rcqxb+CnGXw/dbXhWZ+fMQ1NTOTmvht+cb8kU1
7EE4keixKU08TbBGatkx8jTtApJ8xy33vq8Ech82t+NVSag9vttqofIvyon7hrre
H7wzDC8po3U9e/SoM8v92oViDaz3erGPXxSYdwG8n29d1TZNjxwiauUZe5wUtnPr
0/DkHPn/DwQhuo49AbzZPw==
//pragma protect end_key_block
//pragma protect digest_block
RgONRraHWzkXpxxzQB1I4sG2cMU=
//pragma protect end_digest_block
//pragma protect data_block
P4kzzH4+1e2Osf0EoRSaDthacwSpDedeCbusT/kBoMGlwUWFBslgRsdyzve0oQRe
XTocmwQgnykQBVZ6ZgldDGVX6G8yJAD7kS1XU3Q8iidrh27btMTYPpXYlXS3mHic
z8NKINupQH9uZ4G3tYI1LqMOMTjUMrLfqFw9egBWRxLUrSD8D6TRfbBHxEB3+veT
dozfmSBWykBKcR5vVGpBZIsaalMKm9zJuL1A6k6DyQNtYIXLUhygUVcoLgfYzXVq
7arUaGVeAwHCbOnpbsDTin7mP/rYWYPK2h8wLH5kg9ENrp3IgpE9y9BZgtRQ05Se
8glSjw/49LNb/owqmvXaaXkx37KdnxT1QT5j0VA1YNY1/kL17HTROiK6OknV8zLc
iRdqPIn+OMGcjOpQgcoTOw==
//pragma protect end_data_block
//pragma protect digest_block
sE/HdBm0sQN11wO/Z44swSOoV2I=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype.sv"
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
bAyEGtmk7b1vdVDo4vT9yD5EdZQyFLpzeFjJ/K2SabMiBMyqg88DvWfpgJ7GQi2P
U0zkbKu1gYOYBpcgEfkhOj8oVMONH7wF97SN44RfBvzFJ6ArLUIVhUVz7Ln5jEx7
KGldFwNVdbtG0o5vZHJllMCOdDg2N9UFBgSB7SegCpx0dHLqRCeUXa9K5Val2a+B
ZfMsPaWnuyb9A0HlQ1UEelQqdF0U/rv6MA8ytw9g9iypYk7h6JszIthyKaiowfWB
3NUx2y0IHRbIU4MnZFEsmwgjXbBYaUoP4Mytw/McXenoGJg5d5NnsotMNLtnWvzz
ZF5ux0yW0nCUAZm6sCIM8w==
//pragma protect end_key_block
//pragma protect digest_block
nWYDFScSJReXuOXtfHDuhp6+ZN8=
//pragma protect end_digest_block
//pragma protect data_block
AtltWQgLsEsdvyaGRwk0Ac2v69druaNsUCd7ys1LcaOn+sqqDUeXgLUN1rb19kPF
GLLrPl6P8dQ1wLH51WsBMPIrzQAEL4q+VabcOZqSEsWgBY6LDFHPbi+38Xx0LwFB
2cWm/VylFpP06RN4nRUghOLn4OcMNRAO21+8t9iU7+2Ec+6LAqaFeVr9rhtoH7iH
fhy0ciN6koTtf2Xgz6LGe/ffa0BUAFl0gomFeszFMmqc2Pk20a/BSqwcuRk3q9L5
N/0ugh6D5SQuN/Sl+cb2C/5H2mZ66wbpGGuSQl25VR6mqCIvDHegxke4Z42UlPmm
KfgGMwXLjjZ8KX4PQMG0yiTGwrMqB17bT/FWJi1veDw5iDcrB2RptIGn2SyfgGct
jE0jYVJ+cFttiOyh5yh5Svze5wo8TUGlIAj0UjRS7EPlQpAOBX53N9l07gpFGpkp
cwM+GS18Y0zcyQPUBLLGsV3kEJ9gX6AoGAifjdKKk24WtvxNlXo7uysuB212uoqn
AwHteNQWcFhVVHuHTT6AtvaGZSbR5k2XiWgiw/cSoiZ/wcOH/ilSEh1iC03ulRvW
HHrcHZ4zqNO3zCwfyu5XZaBTN6kfPkrnmELU+Vnxm3kr2rUO6+861rp8U/3a7vVU
77SHjatnk9FElbwK1HnERHXUVj5A8o8fh30nP0IUlm0KwTRquWQIMreWNWVgugPb
V8J+bBHyh52xUxZN+CTjhpylLn6++zuLFMff6QNwKYs1nWWw21I1Mlijv6I67bHu
7RCxuOGrTSSB9vmdLRAQrRg3GDfBDD1c9ObuV4m9ac49iqi3ZuBFGnG6PgcBCI0z
ICvAq29bYSb2NH+XH2s7V+eZmIS4Uj3pod6UjxAf1VPq1NMilQBQqEGcupOL0pz8
d9CMYOtCNm2NdU561I3ZRxlwR0c0xCkSKvzFjaNmw6oOQfEPDGjwsnkjWvSr7/rJ
mHNJ9QBjZXqJZfJGyR9lGReA4fEp+hfQZ0pOp85WO5V7v2LPiyo0DYI7dALdQ7GP
6pgTRXfG0iVfMzNI1VKUzMc662qILQ2duO+76D922eUZ79OgQWCaHPoOcHkNINlf
WUlI4ZM5+RqsvPx9oKqt7Vf2/cuxnSTkd7Z1orExqfZdFzrmZ2hH/gIRFhM2Gl4J
kWE6TdSsMYfBqi141i17ccyl4Ws0j+06y6FjM5r6JQk5dhxCpS78Y4CwLu7p87Ys
xV3F4QJowoEjP4ltco1wbFxB9FdSPoJEq8uhZ0Taz4y4nJgKFVdZ0ATjD8gyTnak
cFtZlKyTZF+XYvnzjXBB/dmOCmhFGhnATEsIOCdOczxbVuIZARb6nNKpPSJKjdye
a6R9pKokzSQtW7wLW5U/dGe2Gp0aK97G+LeKJZ+NfBD96DItfm2ez/KqyMGs3rU9
/5x6S+dF0+EDEtsTJib/gjG8m6Q8toBQ/JsYdg7p1Cat4FcjDYU0/tbDfBPWwb59
hhPX3Mqr1Y7fgZMxMF5FANKR3UazqLxQxRf2Cagteh+XzCnvn+ysPDZYfjV010Xg
JnauhX9lVjqI9B3Id3br3PF4vNfcy1U2Zd/IRIIR8LUaCBQXjDDgiJkihrUp94oX
TNL5NSnN+Cm3mM5owLA+2i1h9j+jt9ym9i8isj6Askvbtcn+qD6hfHXgntCBhvfb
frc5VSQHQT+fBeU5EUjun2a6JzDu9RtYCyIS2H/ZcRE6WNrpcUNUo1DAZi2HTVot
jhq7x5mVKP4Cbr+u/6wD9eEK3YiN2ddQ4itoLdmPpiwbUMhdassgYZu4oD9iZ/Pv
pnAUkiye5UcrBE7M+wTnKlAjQqbkjlAPQAkSGL4cM+hS+Okt5Fh5C8G/CY+uhAyD
m3I5wYWCvSp9MH6FiUjDOzT8SIY/VJX58TWo+oepOux8iAW7xjy7eDNBUkqQdeLZ
Uw5kuKC6ODkID2pjbOU3Kkci+dkdliCiVp66WxNLCzolBcc/KnzsjY5Tblj/Rslk
1FzruBYQd61wmVtQ7geIocJXhak1cy2IUIE2yB9zDBX7M+irtjn/73OID17wYEll
FxoJWjp6dlSKvc66JhLk3t58iCBQ3hYZKrSjA3baej34SI+Te4rEv6JkQVjrhLGZ
zg/x83ThkT0N98K+VD5xe/wmqkf+xlUCFeukKms3oNpGM0HvZBDFfigf+mkKV9QO
A3e968hYPFIxu5QsXAtEFt5d+9rEzEGDPvdVD5OLvRghDYL02WROFjBpgRDs2a53
nwqJx/U7Nc/tbasNgUHd8eg8C62RmZAJ3PiK0discw0wiiGAhfeSKYAW8EJ1wYsD
RDandrF3EvfLq/9GHyeQvyW4QOdGbKRCechaAUq7j2sG7ND2Yz4QDhciSi/jPxcp
Or5YR0fIc1czAxwnFBZepVptXNis3UK0EQ3ktDEN7HS+2XhoOB5rqh6qrZ2P8BNw
TIYSp8zmVQpbAIqjQireMXcRX9HVVwOP//P77sJ7TGdy09FDdR7qxR98sThmc4UH
qXbucrn4+hCXu8e3kdg4EKCUyxjwXYSS0KVTAba4mSy9C6EKD7V9OINoVYCDg7sU
Xhdad1s9KaVq9683XQ8s0+VCMOkRx1iAWAdSnuiL3WAquqO1iorvR5P6vV0TU2it
X33r87yWzbkUH7B2+tPXPPnETr41VcMARBD24DIGOfx3BVrOd41s3YPt2HaTruhT
lWy0DsUkLE4iom8Szh0pW8YRHxc1nod52J5VzPSnBwRWk8CIYKAmGvmrHOSKndd0
kEhw1VEhz4ZPeFx1x7DxyXJS3Jsio4ZzxhcwXK6d94EXXIZaUzdlvaQU+OR8r/VB
0TqHbB0CAqVI7a5erECXzzWKUHKNcw6xy8ZlXD3EDuOS7m17vMOGXO7Nw9LA22uk
PzhuxPzZfNX8Dm2upKwX72PjjoVDv1GsKAsMp9yHfv5/1hLLbhtRvuT7DlUaldFh
nOW378TTSnNMsYzFOJDoF2vN2hrOkyE7WPKWdu22IuZMgkeh6dh35Z81/PYtVyP1
zQt/ea51zmrK7Q41vOcBdsXr61/9uvl9E2ZjMARpgQET77JrAaQcIYHGaKTPxrxR
9SVjc44dKVz/sKtwm0QrIghR1RIe72SvTaM+2z5T/rD21Cw4x7EPQ/8uCIMALqCn
f4fxkEEsucx7FDeY71PX6Z7v9JO1N8y1j2vBC4BWqwncuEF+uXH6GJ+Iv4AY6Q3H
q9fbFcBzquPvTgC+MLr+DcF022LufLwsrzNypPCGd+UpqZVdv+PRMaemslasczZa
KewmQ0h4LDmDNbUU0T8afAc6yRNsfRcJ+pI/VVoqgR8mnj86L+WAgyGBdO61XMXo
Rt/8mUsht4kZsChmyt1mEfNTeIlPgdytC7PFl/qBdsIzegJercvwLzz0SVyc33cN
bx9YWJoUQB7jfxFlfPZi2xY3hG5h4scEU3N38O414+CfHnpsiTATTcKPXJoKwdSu
UHzVAK95gO8d/2Ooyhqrmtz8xxMfJ3jDI4agHGGU7fFerpGCX+p8LGrs9GxgYYnz
MyXuD9mRhgKj3jwsGymDRZ/e5E9866br29ddlRxvdv2/VzsQzR5Bar0dRdRZHaYr
aSNBCs5LmAnfCBfKCWSjZlQ84UVXsSOua+FxTuNruRaW9Vf+2+cJCEHYBRtc6vLg
oUba7WSsnyE09oIfby1rbj0qjr6avZgP3ivDCO61XfVVXuvylk5rqdZWlLXqBnAj
yGB02dZrgKUOSfab0hCrb9jMTWHXheQowDI4ziJoU72WPzjmE5MNoEdoq8QA2XfJ
vLzUsfhxHnsyQ8FdIHofFJt8qahxhVgGSPFC+AVOUraDGUPRUZVZ1diuBcc5YuS0
UicTwkc7/CFaOvGDmKvEXSRxBgEfnN4NgvKbX8RW8Gz2ggUmNHvyX9K0K9oL2IBd
E0BJEbBvLWwhS5wr8poU8o8jaB/d7DKOQkAxEPDYw7USmNS4Xmt6FxuVQ0FFfqj+
eqpYa+7E6c8J0JucdGyQV3omRXZ1njlyT7xLwQOOdX+2OqusMo8Ka4usRNnuDInJ
ELW6ds/Opu3OK2ynDmhnM9c8PcS0WZCsx6aEtKZSoeEK4/kYAyV9wNL/lzonCmKP
q3/vGs3gJrT3NTf3/IggXsNgT4DmhDjVyH13dUeiiNdmTxNKnsVngtPphyjeUM1l
KkbFyguTc0/8BkwWviV6tqYF0N0fru0jedkS1guHa7fKxK/fHSKUgI09B+EgG1Ca
KsADEndvMr7h9/hofEwAdqCX5d7myCrmNcsA+CNz2CMDnB4saZT6+kBUf9vzPa33
vqv8Atx1OH863R0Yhucbet8otIYxkJNzUs4BNE/1SQMHbLzXENhx2VT+5CglmUEI
tPifYwMV9lTEMSukkTAQgkP5t9i9K0+ZdIukYtokAOjv+9Vwaalq0KYXrDWlQCz6
NCkEPSEEZ8tLwRYORDzf/rkOjLfLdVYeWsMDIL6ojVLPd8QEY2rnLo4HBlpvdAuo
gAnPvh7+DHcbSAJwLr3T+iQ7IJ56R/mFwk3lzjW+5/fjGpfRet4rVeYczGYJTBhN
6aTgosuNNXN3kMyEp4cqGXyPXfPBGLqawEJzxIpj4og1NkrWPINCLkvo7WkCZu0R
6OmrIF4/hfUpxkGc7PVM/q/2ys+EQDYk71423lk3ER9QI8+5uiiS99GHJc+MUX1k
5Y7kN+x/5rXnZkiLhM1IccUPRm3/+AEpDyxjoc6Tln5GsP9NLlyXDlmbteVsyUVo
7aZR7CzFT4doP1q6ONmh2b9K1fkjwIfZUaugunaWkRGPye6yr+reDnTruRdkuUCw
qFat7OKAOVBOQHp6pO5GxXHmjb+63qsUtfFUWoNz5YBNAs2oAfpx7T4sVBVFJlTU
EOr4RvfMV9y4THgEAKJhbDc5ojT9y17b2CpL2zGW6H6WDp0RHiPV0P9qI2VT2TDW
F3SEdNE6Zri0qfnSGMyZBOOxH7CtClHL8mShMMiu32a6skAcsy6dzmDBWnwRDMPm
PQ+Caodx2KSV6x1tHCkav/qwLuwGXZQdsGqE11nbRMLwocR+rOpQMUyIkrkGvsH2
m/6tu/ZktIFbJqF/5QsbNr/eIkQrA2AHfrq6cjSfx2n7INEQWjt2FlDsGjj+xhb5
Gd9oWOnC6ZDhm4l82ROqX4VGtaPde7F1K2qHycERuvc16IcwVYRhFEw3EaVA1LLc
9Pfd4etAJ94BVteRHMUi7PBjvqGPqxRSiflqVPqccUYuA51+VIbdsHgrEqBBQyo8
dmyPBJc287MVvpoVbTBYYgSsIj6v4VXCmVxUH2wuF3WxfTfM378YnLyXMmHmuhOK
0Zr8qAnYE8NcjnPPrhs7CJ3oPZE64QRX7UhKv8WNih+FkCMo/qhHQbkr/vHZrXgX
vjS3uxO0r0unR4ermXcqJiNdD9d8g5CxWNU+x0Arn+tv7asbkQ+eHxDigB7Efir6
o8wlUfCZQ6S7yaxkeeZnZ8h1j7uyg+5imq/oPUKMAYU9v48VgqkvUHA3ZO/ZvgMf
Se/+l5VUYZX4fZiJhKrMIj0nFmRjiltiwcySDjRg84pK27FQsQZL0/r7JYdiatd/
s9Xy63dXgzJaTex3gUwCgnFeGYDihOKna9pGuvBKcnqWLZVAG9nCTup7yTnrhBmj
1OwepZe22yjZndvjF5El5zza6hflFaZ2bnWb4YKDQKiOYchYlrioib3UEiRIAsMU
t0aUepdReg8vSfZOUi3ZRhM8FQIzLQNuZ9f2yMQTgM4ylmxA0bqOBK8CzwoeNEug
qkWxbp/L/ij8fO3Oq5drC4Zy0fOeqGVvl2Eh9OP54ZUd2/r+b3/HaS0owtJPy9PI
1sQUe4z6FG7jk3eym90uVZFnBpABHxjjpavzzljxj0424JIKqLLhbo/D0mmasRds
Tt8eUUXwqZr5ml8cypAPLkcg4rMNh4YXdH4ltlZnR4uSe5WMg6MIiw1/CfnMtqOV
q65f0wOo5ig93z39NW0jOlH5X9rBR35O8eY3ktnvnKZ2R/tZYr56ELRjk2gGzx3a
ARRnTMvLqfqKUhb7jVboTJbEYDjqR9QvUhAsdireAll2YvykKtoY6EOkjJaISLZF
gp/izmilbR/GjJxxp33VaE6EnC5GC4CdSezoExoZmHjs6W9yXG4ht2t52PW2Vd/s
3IFxGuPU/sydg9Fj4VhzJn8cNt1RpFQwcFrseIP8t5Fku+j48BPFc7XnDAykB7lm
Q5wX4zcc4XDLwnx8DH9vS6njFYvbceT8Q0U0CLJ7vaCHGZAuo/dsY9UwhOi77KV0
4y1GsqppedeL4rrqqvYwxCHRQwZQ+dXdgl/LvmuWi+Cx7UWszIqy660SEC4W/ZXT
xY6wu0jNgKnx0qobUmMoN0vQ5ncS/C0ZpM9OwAnrBPn4wMgoLjMbVkkmE3fTOQYz
Z9pZs+Iida8IGVnlCutR3EIvbSzimSkOK9Iuby0uMs0JmgIfXf324nQnY3jptVSr
jucaOWbHRRsqJ1AZjNmHYNMGsgyq9GH/8ThzdhYZZ7f+rL5cVrizw5YVpZrVoZ9r
M89aINubpQXqBq91OzoUWP+c7MB3IoO8DJzaor5MdJWcwTQI75h3OiKQChD/UxSb
OU1M1AtlNH7kOMWXI9nePRmk8MHoxh0SxS++861WV5r6bFH9OKyXw5wCG3xBILKG
5G/VXarhOKSl1gGT0yYx0MtQZ6n1gmMAR4JnDW5ADIU9h3+3eNhl46XaXqoDwZFD
u4DRhcsZMqm2k4GollcsVkYIV3DHk7jzxXfaJBwWV6Y6dFsf40JZbvGvUTvbPc+e
vCNxbw6ToB38HpoyZ6uv/1TCnHH4QSp0WM0VbqCJQpi1ElXIjKw0/oexNpdRKYQk
Gzbq3PtHrC+Lmi9OTuqFGE+HHjL3wRwt+1YbMAQ9Q49xEr2VLuHzG6miW/8NgoH/
F0uaU76T7dG7euqEjMsCJ6+FWXmRtmz3rylYuJKhhSYNcIluJwnTC8rL10JSFNz/
yqkwf25HKymMPqA3cf/D7nBdLXEVEo1CyRmliBH7UgNd14wM14JzowEMo5d68GF7
LKOqxr4PwyBXbvvn16xleJ5b1L8+oa/Iu8yDFtl5A5rLf2gcDe658H+zP1XUA0tr
AnVwRC8EvacxzXGK21nSqGLAWkXa/GABgm3mwukX/9Cs0MpC0ilhCf/ZNT0PfLlR
eciJh1HtwPbNvdF1PR0Z/htpU2nk9StIP96Ix3CbVSGH41XxJ+oNsYZyaEgYf4yQ
I+9daDLx5P0v0NlL4keMvB7AeXBa3uQlzgKjKuxbxejWXI8n/HLHtkGlOSSd1sMM
3P8MpDVOUgnuGfdPh/uL2L+XU9tSyf07pLNYpQqOSI1kPOQL9L/TV3Mh8euAH4pp
6Ovn7PiVx+/0MO012flfDYgu/l0998VGW0WN1mBhioE4FrQDNaNVAWWiZqhjvrrO
8JT+0PwmDGIzVqRpOUmMB7ykxzxNz74agr+SMA45akHm/GukTm0dV95tGk+NR8VA
iwu6EiKMR6VuoZ2Zhd5Bei/G0DpUlgPlUVPPq0bIiJi1GfN1D5jhFdbfsmsXeS6E
xOrD63LwDmktueA8Nyz9o9J+J6dMQXBZZugjZUybEHiJrxZ93meeUqAo+FA3Jx2z
izeAhME57ygvcP06KUfbS6giW4CQAUT+JpOVPYdC6/BOS8C/1vBSj3K1kb0crXZg
KDEeLv/LfN4BxBiY64efCZbveQAiGIWlgVip3IM2y5JiejaTsFS3ImnV6xr0HsHH
RljbQiDDjTzRNxzJwFTbEp10H4scTQqqvYzKyeDTZQHIAGOEAwqAYboIZE2FMuQ6
jINzGh9brw2T6kDEO3Isqbf9tACcmBHPiHnvlpXW3jLXktYsycpdMBmhWg9nLWY7
I3+pVqv2HefwpyPsIl0AB4BePhKSdpG12xpC0AJNyuPsVFcUZnaZnbYHiZTDF2zZ
KjG9emz+8R1InOk+lGBrgy710Xm5U1CoxKXGYjhWl0YYL4V0Ny5/wz3l7lNEvjAa
8aPh5/RuryIjMLxJzB99TLDK2s9JDe2D206hLMZfaT1aZvBlg20AalpNSwTYlsK8
3z0fkEEIe3uxWjyUSh28PV3EkaNY8zU3b9vFnjsi65ZdYF/bPcpVlLBMRdFTRifE
Te0f2gTyezudn+gTxgoRpyCYf/MAFtYk1oMfoXwEccsf7bD0BQJKn/rgBTNlD9ax
n41RaYGM5cDzg5dICdxaRt7fQB9ndsXUfOVHnsPo11ihwt5o145Yc4nwMcnNrXSN
XROp+zaTa1OPUu6AQURvkBGkal7wS7acqQCRB/O52EKxlZdfdgH+4hQMd5MigE0N
EJDv8jA20BFU8vYsoijQlX4CaSbMQjea9Mnb6R8eyq4uscjsE9sEyKGb5df9kogY
SEWn2Swye8NvWhj6wS/qStSzZJu8KBHlHqulM1V0kRzb3ADDsczeKwbQSIwjXd41
vo/6bsD94LlI3Ru3rbz2pszz6VvB/J2e/yxZsV61GgwkHAu7WAXXPt7cJMeXy0Kh
5GY6O/yAi16rvbLp6JlyFwo8yahmWCfKMX9qFB+z+iDJoil5kpYjkxlyW12yPBUj
33cdurFR24S1rDbOeAsBX8sZ1TAnnvQ5wy/L5iVv4UgFzNftpHFWB48PWppdLNwn
TEescqAeXJPUS1Cng2jiPZwi4Mj1P03KRcXtB+vPWTxtTcQ/V9gV3lWwQWD2VO6d
CSRIcHGAt4sh5WOBYDhK5zgFl5386/7OYXYO4SzYZwr0zK/m85CeJInZeE1xibAz
febsDLqt4y2HkkXmn/LtUz0dyaGTYZYgp6bNOBbA8ZI2mMrLKqLBBdhQFPT9h/Qg
F61VrioPrWRXV2rGKcNuJQZU+ZCGZ3jsw+bh/XVpHyFvRdgy94Y5ln9e+onbsZxR
RsHChxE/BhtXm/vQrPpyP4DQpcD7O5xB2dw1+rPsL/dYOCa7Ziyl6mHBh+6QKaQC
MDdoIEFTXdk0NJ+QtikkAlD2Tv2lebpfzz8Juiis23uH9Pae1Q6PE6/cZtf+X2Sy
SOUvpOEXwic3EXVXS8x3zFmS0Td8fWFvs4SJ5xzZSPm2rHoQny32LYecbKn7G1Rv
evdOStVBZ2IxqFxcPg5/+axlYoQg683rFiF4vbRoVFxpyAr83xtBo9FsDXScF14G
yTcl3snyIhDgl3T0qwuu0gp3CfBQ51n60JSaKOG7UJxcat50ejatZT09N/vtVOGu
rr4+xITMKDE87Q1BENE79EZgTaJueA1rPhBwdezbNCtrwA51I0q0YvDi2Krr/uOk
GgJ1KDrpnLny+LW+bWXFRCaGV2X8B7qS0mrZXbbSJ0MSDek1rxca270Mtf3RaEgK
3E/ttQap8vgS2Wdu+8cc/mQbW/KpX4n1ggOqaUubKGLaQvnh7Y4JBIMp/3jVX87f
iXmkIc1D0ACbdXWMDuTFWGMVOVZTK56h3m2tZQ2XQgzgfrRlOf438hOeMLh0Phie
lYMISUp4tc4zp2aQO7XcyBQ5F9oEoEBkGynsSOEpr4t/Lh/AiqdGf2GYZS0BUPwK
SbhCF2+a+C3BlyDBUUKB4x8UPSIguZv2WCxdmlF5LCBdt/dNtmfTVP6ss3tku9XL
NyO1q2dYTOIJgQFtQae2kI5BzhsBkx7/S6LnSKnxm1F0bLbca5I0D8fF4eMsFosw
CnNSe5WXyyzdw6eE6wIiQX5iGhszN5cH7cD62CQKMqC4J9opTvt3kbB7cMsXJ/LG
NwLgdh8XXXB2erSOAIODCndFCKgQvWSpt38PvQyEtwsapbedYsvltB+Y0Updbkki
+HGm5Y0LKShi7OIFKInBOVGeVfF/42TLVGOeNMlrHHLJTfcHlGVDMkIc+/QG1XUi
PRBZPN8DFHT4jI18mv8AR/MssBceIhWOQYDNZTU6hBjC2bNmpop4afCE8qbpdxBL
0ixwsd8DHpVv1GiefvD7WptORjcjqkh98AtlsiUQ3O+y25sE+2jBzBiOyz4gy2Nt
5pGLANf39GVaRq3BYJOY00+5p2LUk26o5aJVEld3C7JnivmLkOyv4GynBF1UhiDn
rREtgHYGdqkq+fRX+OMygl8/YUaYz6mLRLcKUFqF1db+CXLw0ULVuFSNU7SW+BaZ
vmWQbYWBK3C9CRMzOQp7j16hfPvE96ki4dhW9VX5VmDVMhR5NRLYZYjpyFs1qEhB
aNbQPRlQwunKEGEqQme2O+Qwu50djEGrJRW1XmUyv/DriIOxILjWlFi4btUob2jX
njeKAcOsuX9cUbf94RYBe9vUVlVvueTj7i0l5ra1NlZZjmwWdnjn/ZYmAMCCFROO
PrmsJxkzSw9YnZe6NGWJYLTMyriJy3YmDFBk51TBzqt/YpyRmTFtuqE1e7JfQrBu
9t3ONMcZiNyW52uaVYl/970w/7bGq841StsrYVNW7yiId3H7CIL8NGPuRmvZ0ub1
h6niQSsR/NWE/mb8zkGv6VXy4BmhhQDqkONb0if8OHySzhce0xzbEDWfFRD3K5Yl
oH1v+rOcjteIYpZyTNxgtnW7jGiZ+U6wYNLFIBh6gkBIWA8i2SjNFT0u/m3isvaf
b+1eq21QE79J0yIV2hFf9AlngbH89pCbkRY9Es/jhvqeNBIRfDOdTFVf1MLzoPek
wQk/THDVzUdazIgteyHukr9EP7Bt4iKGf4W/o1oxeXMUmNc4fWUh2mId/hRFW1AU
YvHI91Up3P9wLmlSONGEKdQ+syuf1rdWoCU0VZCWw6SlFFLA6hUv6ULsSuLO3eN+
b0n8AoghG23MZjBpLCYpWumxFS+bh3coKcdvRUgH1Y0PMHIFRmszSIMrgrGMtZB+
JjhHJ/+V4MDzcrTnM4DmZDOnk8hjXNGgN7/UU+vTnNMBgbx4HINkJesGG2ltNKxT
eaiIisF0BKttEkk9QcoecwqWGu5e1YRZ7lspaRLrvfAJiXoiugQYuk/VBkqF3K4V
7YRkySMd/oMytTmjrKk8lRp1UShNgomCOup2I/j4aHqAAsmdOsrUtRiGOE0UM0eB
xbq0jM/iHd44gyk/PW4nADYTZQSyHIwCSTbK39Z3RdzuVIPBfQGLG+gJHMKMAB5W
p8lehZYbNnwf7e92KP0dHfcTR0D8Fb2yLOBDMOASngTJTS7XyhOWJgt8ZyDS9Zd7
cP3UYNjB1dvkCUNBr4ElQ5bu0QljDBSkZPkN75Sv+GfpBTEU3WChvAkcJg7SUR5W
mu4RzpmBsqNhJZpHl/sRTtyENdUJctgp6fZn3E5/8mgZKxsT+t63LMxB1DbZUSz7
xMrKgREbjhFxjv9MpzAE5cfevBlgKksyfQao066TZJ151NlhCjM2uedMvRJTQOIl
oQSBSRQou+05Sf8XHeIcwwVyBPFWDpnn1s7fx4oGCAMqpVYuP9DeMJ5UNRRS1c0K
VpiOjYLFlfX4a8jDvjuIC7GfS51mK5J8Elew2IndmC3ZDC4NtnqYho/yTnb0md+v
rYBZ+FT7ek4TVyT08hDDiGI+WdiBfU1YiL9f/3joH6k75ylvPTgwzgeKBiMwmdD7
MUid7e88e+dPzvmXF9ooMLPdWBLvallNMH2hO7EaT1PLNs7xYoXVQrArvC4JBO4u
WbhjpyXPcm1Ipf17VqmU7Qgpp7Ezxyzn6ns3nqzwksSXkcwI99gyg2ZbAvtlg6Kc
1whcwuKyiqCvXSaa4/CWcIiZmoLtxkOs6VWdUQT/zzrxHn9WRSy0OEQUa+gPbcjq
PlDEDAsa7rgm4eMPHa3ftygEFg3gKTh8UtJY3KAKQ9TmVdEwb1gNRacwRtwqklOJ
0QQfaJZobq7T1XfUj/V7BfXCWgWy8X+WTlC7JgsqpC9aRWT5fgYieRl4oDftlqnQ
3//VNDlAx3bD3gIOvcIU7rH5Ur0xYst5wXv0u8L5FKc4vGJ5f6eHMadsjxTGOV2z
DryRJ04g8LnJfkKDGCMqNW3JVI1uAyrjHE8oVpyU85DVQ5wLNPS8bfOiD3vvNxzd
6ApKJf+Ho5JBHSMx2Rp8F2GPppFfZkf6UCQBjf7wnaTje5dfCZTeO6wICilP2bTi
8CACc3j4GLpH9Vq5Vl67tn4hy6texVPxZoZ6qFXy8v65TwzP4CvKSqyd/igJNfjV
a0TP/+C1Jt3whWE/6rwUTMn7dS3kfhjyPGVZObKKvdreXr9LuiioB/jb89Py7Uu2
SpxADzdZ2m9Jmgt2pjUarJKr9Z2wgh4kt5o/ZcZLLE05p1ngOLHfoUFRxFO1OC/+
Jp4cbIHLwa0nwoTu6+npZGrHySU+4DQUGCj/t9lSUVE+uvHcqVQZ6yPE64poV0Rh
V4l6CKZDIbzlPqJbdlW0oWXU82T0m+wmXk1e2TCxmV2S3qn6ySrXL9tjOanZlSjF
MHjy/8k7vFzpHkm8PmTy1Y4wvBRjBkeoV2vmgfXb++Qqr9O5zvEF/27dHAoq8L9j
k7r0DCTf00YtlXqsOvqThymTsRg/GkF5oThUJ+ICv/lLDIAERmxvE7GKNRxQ1ybN
vJ5g/1RQ2smFd+4seSbHwDiEb2jhq/jlL1In+M4RR1gDv1SwT6AUve0TivzZAFmV
Q5ecJIGgmiMbfeQ8InjWF+DdOr2lZLfPvMhwQ3H1nn+4yF+hCY74bLbov0EnxHvD
qCkGgot6wr8bmWSdi9twHIFUNr4Xhcx/Cg3JcXd0OQp1/5jfoC2u9Y+N1C034wDy
GSepj9EwG+xKPnXL4+GOJku57vdIC982e/02sJPZI3/y9+7Om03SpIJawMdd1Vm1
9HQj3v6kfegLmK3Uz0gEZnlpIwwP9fjsK1kLnt/iO03RaLrI8iA7HJ5fahMMyc9t
FTEVxlIhRDw3fMQ44hJ2qgFOuixtAqXPSFMr2332SiGiNeq4NFNq5Og/tKZDM8x2
EytqnT2scieLnpetIzURHTYAS8TNGpp8YimJGbwKaeZtpkTJuVzSdZtTMD+ggNHU
fIqZpsp1AJfwvM4ipKlecbgVEU7V6Olq92D/4ucjcoLYoDlzJAjZA7RDHxpp2+tn
0tmi9ZX5m7XR4yEbUNdrRCHWmkb6ELZa+HwL1K44JZWgHkw93n9LaqYU9bGBnGLM
qriNp12ANDBlMCpMOlqMLNL7c/hmkWrwxOTe41QWxP0z18gYIkZxTyj8z+qmpomC
XWAdMg4sIc0r13OHGC23OtN2w+48P0wu/Z4pSkLSjYPlQvf/6bmg52C1+hKechaV
iUJw4cbLsSV7VuTL816eePuGRAdHPm3bAXxBi1FeqDKrpIhpxOtO8Lx0Jj0TzEbz
m48rjYpexXjEK8XnUMMGIeZnqGikX1+cqsaINcYNQHxj9RWZzNIV73JKPG7gYzqO
cMDl9MCE5Tt1m4TNEpp9CDaIh6YkGztKmohpG8oEmISOJWqBMLLkQJPU6WnrYpSp
wn6MG/GIJZEAkNzr/gmFuCJWVSPxEXVHEgF4rKEdLFXblPXL8ysebFdJyH+SMfOf
Q3rAvqQa7iMbcFvSus25Ffa3tji4BehIgehnlgKJvnYO+ByMxSxBFNxfZilavh53
ZceqEcaqSOXHM1NgF8o+q14PbXcArHpGSzqbS9TWTLHzgCjyCavJEUZQf6Sdqze1
JsdoSdGBa7GaLXupRGLFebcpO+YUu4IIQbOU+19/BAK/Zl2vQAxXeAsEzUXJ8W0r
EiSatf0mRVNqjUezqy6ER3mzilaACbEh4tN3Wn9g8LGrRj7FvdCR37cYx2vUczUR
8RxvZ2i3ar4n0KGn1L0k2/cfpwN8SsM5KHg+dG6U5DgmmjsII+oQOecNXtMqdiQw
IT2yu4wOgfUiX7GKvzFAO9IO24sWnyoXxBuQhj9EgmAtGEpTv9Aa6TBLdeD4/F2c
M97ve4u/k7lgwW+LQYOGGeKL62UnGpyWQgUO0RNdj4N664GOZ7bxZHxSw+Ut/ZPH
n+HDRDA+gCLwoWOukeUTE9/9LEELW/MuUH2VZsZnQPNOVuNy/rfbskmZpBC9af4h
pHRN54GsRqlSvMQobMruJom9AtMKXt5WHiW3d0HnT+kIF48z9LCBn0i4SSVDhVWz
y33L2esAdOpCbqvsP1/QXYdsRzMwxgTGrw0g2nZLwnIWcuW8xpM+kPmGcQE+jTq7
FadK/340q16H5jryHMUbL/htaEJ5+d/mEKdc2u6/0dotzYuLHPJIJPWC+LqAgQM4
arwQwJgFwiDRu8bsO+Z1Uz3vEjIL87dMXVqJ0zfdhCrEp9HXuvnH8HX4sBg5f75l
LrErQCKLtezO7umTACin2K0jT+zQdTMysWuOfIyZ2YiDgN00LN+DI5wb/511+0Jf
fA+E67vKjwTcQPH3I3p42zDM6Fiex0vO3oh9oioicF/xTM52IWAl9O8AcMSBQhU0
BZR3jUUNLXQ9x4D54/Q7Xg/MY/zO5zc9QZDDhs9T52sOHKkvsG83Qnt4iRGAjLmi
Cg5FRjW2jD+ExXznanwV18sl2PAa0HAQ/OMY52f3IgUVXYNyhSsPaOaz3a79ujCr
bvYdzHb7Py+b4CPGOChUElsUwCIBksOMjFOZ9yaOzyVFicZsIMRm9YtPVkdg8QVl
ZQVx3Wv1NfmaYFc+2MXXLOYm6ldyngGT/IFLtrYH7BCH+cp3hn2SVKekvox+YbO/
u4CksB7aQriGrISDjJznuPzAyVIQ8uI84Okdj4MNehPidhCq8SbCVhnpSmwl9lZ6
lkJkUTcl9XIGXeJJyR2NXBrOjCCf2FWganw7eEue3dwSYLRtqxKg0iyXWnSwM8Sg
+s7LVoWWzHXSCl2edqHHtypz6JVLL6Wx4WOywKsdUOD5hTZPKJNk4SQM8Z8fQDOn
Y9TBMWWVrPYqEGYBzRmEN8NM1IUBeVNukAg8yCAlKZr44PDJvQI39UVATNZiBt2A
zio4S7xr/cSL2YTV2udOo1aQPkP59CEhmXSJXt8aKWCBu68c6oATTZlHuAFN8S86
Bwb39xNIJaVZY3KvZFj6SIJWXHKz+9t0fdqPz1exQDx7/PgCeK+yYh+yyfMN7Ec1
PIe5AtUeEVipXVt13dLLOr4bfTZGpvagpRZ2OxJWMNXDPIdLChAIsOqyVDLZBzYu
JhkJ5gXoUOUpSFuFeoEpHE3W3fNLnW/JJKF9Zoh3SaRVWH2L11OTxU1qE7e/QxgE
xe9Nsiv7CgDSbQEO2S9wFmdD285en655rGsPMDDCnoca84tRp2xrJqb8z4XKbMp/
eufmkSZ/eOmi5v925RyICdfSxFlr6BAsOJ0+BmusPk9O2olKomcdhCLzsT4uHLmO
sb7fxeZ9m2EvN06oORn0q4zMrwZg57vXlcji4nJX3L0FWUtMKw+L5B1XFYixhlRF
pXKm6UlBT5mEN9HNd4zfoWMV4ztjiilGoSse0zHLgxEjxkif/50+SF6LQdZqgGAg
x/QuxZbU/xY2unRyktuQyAouHGSOELTlY9ucoIrHNpIkbZCUM+ONtRaw1M/zjAMp
anQv0CSTVNTY2R4hHEz13SiJX9JHpMR309AJ9xwHxm4clUshF/0lPnoqB8Ol98vB
iBUhZY/KUb9xzPBOiFRrr9BCeEPOq4nzG2cbctYUEjk4CIRncj5xopE657vZ8Xmj
0twulLcXTWTNvHRUidtu0poU6i42QHoqFFEZ5dRjE0BIJ6ZKOQdDAkVh4xDLx3fe
lXi78mCX5XLfLxOU1okqhwWIkoUxN7miS1igktJCOus6CMWnVmX/1ASqPJ4dlvm9
8qQh9t7PKWA/7BrAH8NAuW97Rmh60NSysF+B78/ns5LALg/O/rCMkDAJ6yb+mwzw
K/Ybu21L3v2NBmEfA+Vqlfdr2I2FiDINl9pIg3B0fRI8bXs/Web9ReeHHM+8r5yZ
wWSc20zF2vX79K80B5J/taKJ0U5HHqq98Sc7JPyby7DL7sxsxSgxAlMagsPy8Xl+
Q5nmUBkRv9QuOPnS5tGsfNXSytdg8KJHq8JNIckUARs5oUxN6px80U2hxOCM7Noa
QTlSQmObphp2ekLvBRX+ml71CvMXe7q8FabWkYQMxEaBxsb+pf9xNIiyUeLyJgLw
b9CsGWoMttuGjYyYhIc2mBiXtWKWgwA2G0R1MiQESKqlPbpWtuoK3M8HC+IXS8Nq
CycTZpnEWA0xqbzr/YRV+/kWvIOBVcljBJnNPti0M0LrvRdPXwhQQsvCmydB7RM1
G3FK5EmStyPSq+89jJXH7MXgdftQv+lK/2k0TJaet0XciHC8T4QfH3GlKwP9zuwD
IcISIPyNjF6N0cJ+H8rNrYJBhwroWVS8IRaYPpNi9YfzQqTRy0KgDQkKWG3rsxE/
imPou2mTjKHIYToVsqywRHdSFDxIZ80OSvVQudkICJWbUiRwyAoyHwT9LoL+WVJc
jRvKJKBhzg13x4njhqZWVLjHEkYqySS3GbfHuoitXUwNf6v1+auoXRtrwQxca3B5
3mzjOufmWL6gKhGHgA9vU4gQN78gC4pFNZYDXY1OfGHIsi9nyD6cBpbtshdYOgfd
Pcc40vixYbKJ83lwQrYRsIttgLUcr38Jpj8OnMxE1z8D7vtQpF0BXWt4RvW+2VtV
2bS55nrVhfXRXNjyLp0l1p/riw5JItDDRnKfeo7N/4NBChNKdSITGRaXayyLnFLQ
Hm0udwooo/bLyWQskLyuo0Y+5xhXr6ujoFYu6Spybbell+rRdnPIRm2C+wSC8ydx
Ws093TelZRkpqs0VcPwwVhYUHCHRqSW0tXZ7A7S/vr6XqeF9uYTjPBzQuME4SJlp
tdG99EU8qIDAZEHNG1OO7pvhEUTaiG3Jye9A56GEr2qF/gybss/7UKl6fNZZdGgt
RwardPTdKqO5eABkjyaaWYMmv1TmmjOUDI1ndRD+J7zP/uLvTctfgr3CCC10pXUB
NRc+kUiDuM51zhu/V4O57bvvZsPHTAmKW3J4HsZckj7i2n+DiSD9AsE1c2J1i/P1
y0hz3lBC8mFijRy+EDgFETG6dxeXl4gr3Bkwq5fB4XqTSJmJoRzDnnrLisicL0mr
mR+MHBynTBxaoVIsIiE9KXUNv+NTcoerEo+kZvz7kE50LGgMBSA/T/IzOGOdcw5A
n/P7VlDr7SLEheHkgufdzwIoDP0i0Amag2wg40lBhcIiKmDfqnbxIlcFAPL2pa3B
GbwcwcbKL27MjzNuhnXlJLuG+Ayj4lJqc5iT+82YLfyxAfYWh1daFhiSo0bfPoYl
Szw+xgQPdpn8MA42lwDnfFso1dVKwHMmf9CWaED1NJpAv77sfINNUtE6GBYL57Lh
LM+PGeNSg8Xd/ThtNGPFAkrW2KURfbCNyh6BxSn1++IxEJscfHDWRnOf24uex4EA
vhSdyw0TeutEFmyH7OvkJGQ2gQa5o4D4PzP+u9XCQQmORUfKvANM88nXpmsooxoc
BlV8lq2IjJjTm63Sjy6RKPxF59ZwRExwCiVrf7w88GL0JGF1Np2yX/7WZM+OqHY9
sfaBr9VrdMJYcCrJE/9cSL/0uISyGM5RDD1rZUtnzUFCxYToBrBZR2pcxxuC0IzH
dooA+PV10oNRf1nBrbIuxkmfnREalVRYxsqDdD1dWNSc8i3/cPwl3LqCmOZwnE1p
n0eR0mopvAvwXq2dVmxF5v33SgNIxqgtkeSZDueEAyUYC53YxE7g/JnjQsm4eKpt
z1uJGUCqnJQxQ41AhTWnDc5UEKWWAvEcMBTj0fkKl0m6NavHsbZwaEzouFWSZ4uW
rGJ+DnY7ilkAjGpAIuktSDhJ8wGuraoVBV7uFu2AB0KjmC63jRzl8gRasNGO0AvX
DfPbG55nEao7+m5/ElenREgrJT3JRcVMDYlc2BEaNZc2OMF2vxI1j0Fp94M6zPV0
6KVN3i3wzqEqwFGVscVDr1uyJbLqhLCqvacyNgK7a1+VrHAvXPxNd0r6FHOjBgz3
AMS3YVoFP2f2k8+wP71jbNO8yPjSa+r1uYgYWw9lkWwhQG8TpXiD8KmD1t6KttPQ
gmmzeZb8eqdlhZN8xwtDSVtaCD5DN+EyhZlQPmX+N5x2uaT10EjQ0XCsfL0VZP8F
GujbuDjV2gh8UPutpmjMLQz5KQUIpMDZMZ4XsLfHU9A2yuwqPaMKBsCYMeJ4z4Yx
dMs9khFeGfooolnvq0+luzbgj7Mt+Fj6ZljczevMty85vtYbNMMG129S1pS7ERLQ
KuXBPWptMKyfpf08ByuDNG84ApOIdJop7SO/ShHNU1l2O47om/LcPwPzvHeAh//X
hJJ6cZJPELJ0tM8sGl4odQyLQsw4/clXV1SOxOX5cyTDGRg+W+48VJfARppWe3Sc
KtqkImkBxVnm7RNleEnBiaanlAAcTqtmGfq45apAMCC+CX5WwOtZogsuX9+QJ8WD
6rRDdqPCJPiFGP8+Np8p/V3V8P4aUq8o+Bx4pC9u6Dr/597m4h/mNY8kyhyNgL4R
f6dTR5PeReLztlCmZer+q4oIX8MAUYcTexWZCGoyTKjQGlQu6iEwhoDJLhOS0NF5
COqFupZJX6F0pupV5cEmm0xrd709v4VoNzv8gVg9SC3Eq8/hrPD6f3BG7L9rZpkZ
8ICx7lroCAmQvOTzMIXOaXzXTZDvRPIPbhdesB6sRMTYJdzNzUBMEmPHaXBgTcSC
gcphN8NvNrxo38A/VDFzoBcgxZ48ErmQHfCOoy7bwdG6bMA4dww0PFB5TYeSCkb2
XZfz9IZzpyb4GqyvauraWjQcmZZUWT9hONRe707HxqSTUK2Vn1DNygAmA7ZTGJNS
CmuN9Rd9K/JqjWNHZS7UrRS0nMeg8Vb9a7H2Cngm4SBzoUBWSPxezX4qMaEw03Eb
MShFwCOx5HuAhSs6eVHOCtEYNfDHJIUOWFhdkC7hJjvBBHSERoRkMc+MGm/nRqHV
eXKZySIiUlw/aZkXWXVRKXt5+1ADcRC5i8jor0Xo0UNYE+k3/QxGp18QKZzcqexE
2SBZb8xUJ5PQS9sYPO1Ga6PiJh/luTwXNBStMwq1M3m9uwSu9eBtGpXhMvtoGJ4p
isxu1BfBiIR7Xg5wAHDJe2QTrRbWy9M4E/GzmwScBo8aD1qHNX9qtUYZSGhtEByM
zvBTCT12riw+QLs7fN566gjG+rlnfBi4sklZFV0KbE/6aSGQ18F9d6r+A8bm1UF9
Sm/GM46KWPPlDMOmNIM9S2HzftyBp96Bk/6vOp0YeX2QNv1CEbRq+Vh+2NoJQV+F
OdA7xkXGqLZVaf3A6xXZk4K3Pf2auriuNFVc68hpVCHnyNZz1hjbpf3MKcTrWf0D
uALWG/37apZdKtm1/jeo4vve7TUFyokr+G1f+g9Qy/Tt4VM9FZel7p6e+DIVEzvC
Ty8GCgOFT9zbutASaFUPT6jPQDRP25IG61ja1EUAH7tvk6WogGLdTRGyodTekSTv
2/ZeAKDIzDX8GAZp7jmPyrqvfjB0pL7Ncyob9Y5u8fVSm//E3h7yM9uS/ewveDnl
01g0i2ncqhjdxCru2Sh1D8sEtsh2PMkxBkhalEsd3xzLieC9ppxq07iqVsYlqW3T
UusPUxAv8heaThdMdtrI7h2tfn18PjsHP/UTnluah2hsmEwGJULTDwJw9irF7uOt
nSKBbgzA0MHnTj7ihMrIRTOzndoU/+hE+fPA3yo9DIIwAlLlz6gk1TzeyUiDTTnS
SfdhKwel3xGEdRQ2V17ss9QNBihbbUEVUK595G51i8mDKh5xbNf6ttseTv5yMHi4
TotvhSATHSNOD6ihNntYPcU4cljxpyXvRcLrN7jBPzJAbNSLTlKlWAHMt2PtvIX8
2umJT+5gUT4Quz1GXcV+PngJJdBOc6jfo3iNQlKIn7zA8oWd3m3JUwBy4RFEqw69
nDpA7oQZ150AuvKOIrsqK2BO0+Lm+bEbXrNI7oskR3RO0lrJAzZ8k31MIuB4w/Lm
oxCaT8VgTf8Fdy56E5sb8G6/RNlhK7wMLYn/TwTS9b67OH0b2WPqbxaMqbfC56M/
bUagX1FihPhbHPXr3EF7cfXZDVQ3nTeQRp6nFFWfowkXZsqXJCciXXr/jJWjZ92F
qofE9gtmnJ7v9B+csKCITmJ4SdFN36RXI8BHXk+MRAFBXsJDgr7QpQi9VUGpkoiO
xiEeZOpNk8aeiQ3SQT9ISutmJGvMBr3WAOP5xtqnn2KaoLaXLP2ECLfwnHx0+1aJ
tuaxrJynXojJqVOf9fQVwEeOfnKqRY5ufVFZbuGkzgM5kWlDe++yEQHui7RMiCmM
zE4BkVjR6RNqQtkvMy2jfqjB+P+ghsuRBLj8ERdUkUN0jh56BKdt6ZraUDEFbEW5
Zoq4vj96/gqcjjl+uTTeCkEwYkQrkBpLK0Eoj7BUcqr+MQO4IAgJgVwQ+a4gvmOB
Yg7gfiRYMXRY6yQpJCi2xWaZaLwFHPab7/6llZumFkq6PLrJ5c01EsMCvI96YEWz
+jEFV8XnZxGeDThJ0hvLgbfMcDn8hAZLs7oYlL+oIsyjibN5S/td4NLWmNrf7qOI
EgVCiNtv95IJOup//TpProUwhZf5Luv3hOsS5WptTyWRh2D+DvoexbZUHn8j7I2r
OX8qoF0J2EA+AQu4FHoSNoZ4iZ3jrvWOTZF8bduC4dZBio1NtEDcjIqzn0V1wciC
2fgFagjUnKtKasB3GOj6AqXvWyrpIlmA5/uuSqDj7akUPEH0H7ntIykuyOsqbVWs
VCF+QUbHCSjcEStilLATeWW5TpefF4nRhzS2AL6MbrZRCiTcBVGEy/NMurfST04s
lE0HNusVRSqbQeNdfphRkgBZFW9Ozr47Ue7WBzFx5NxzVrNpeO9rrtbr0H/cRsyP
imEjMCGKfaOdkY7X9ZuP417eV98NXen8zsJbxFRP+xLtCr9g2Dk9RHXWeCgvjG5w
fXqVGPcCpqVGhYHK6PIapTY1/l8DP8O6+lY5CQnVspl14w2457EgC6gOFtSGBFnI
TqG2L9CPECmlIerZPoYqwbD/lM1sFk4pYA+XTUyG4k/3IC+6sA/Xdmp2Nn06rM+Y
VKTYnmshOELaRzt1VQ5pz9zAgoO8t9fxVG5vWG2pk31nXOVLPuLXMxK6NPJADw5b
QtoV2Ym6u+3KRczxiFjoOTDiKcP3nKWA3eb4Pn4L4GJJTJ8WdSFCs7AzzdEVTJFS
lEXFcIhtnQ4GHIaIlbyaXancfKOlZ1n38shKIgwx6WZ/y5BUnu+QGs6DOSKuQc59
9EenFlLm7cHXbhdCVu9cNVM01Oxp9YJtNNbAEEn+05pu27E9np6AoKBUlorln4Da
A9zq8FafkPxlCRlKH2ksiG52XHQ/MgAszYpxsRMDwQoTAwiCApSqnc7zN7V3fnik
oaQPQj2xlSlTTRC0Ct/MTbYref/b7yw4VxRRYFHKNxaOCxYQHL988jfQrG53/ClX
uHxT82yzYUvnZgfbgzZOuhid4KVO0AYaGV+zCFzST1pRpKATYdDSCABI1oCRL2Yp
UUS8HKpOGupKxDZivQiN7ZKg3IGMUcPMXxJWucwYg/X/aqOqXQrkfl/W40GE70TW
/w7PF8M6w/kb4v1nXE6Mu7oRGpYwTqVc0y596Dv15KZ0/tvZY/fiFSp4iJgwNPmd
xwqqziwU3S1A+QvcpBMpmdVrIOY4EcB5HLDqqUVwX0k7MoxRZ35QlBgp/DAhXDmi
uwGQWJDJG7UCMEVpA53Il4o/4WYNbt3QIrO1DO8GXzR6ldin8RZ9ElDzi4xzbDLu
5dEubpd0+MflBUjo4rYuyxS0rcPNrlRXPBLLukKPekr9vClwYCpayMJE3dCojwLy
gsbGUwXZaSvQ4j16dh6jp7WJsFFQ1AQShBQALjAhSD+QbnwkREdvLwHpSYpVVGg1
dBir6fnzbnZj6sZEYA8VOWv06f/mpVBb5DBaUTLc1g1MAylkwnCwdS/4BKqxFfST
qMhpaSPo6kYoVc/UCRMguRBgpsHBa+6QF1moMuIh3uPZqMQIZ5nI4Oo5GpVTiO+P
+21yz7hz4sNegbrynYB42y7pokiJ+kT1LWmDb9mwfUeHHFLV4KCWWq7QEZ8fBf4M
D3yu8WtcnrLnktEDRsjk0VqzRy4VHLD0RGuVkEpkTHin91le9aeUT2hIcECDMvXL
p74fyGsqG3J9HxvQPg+uThgg4y2MrJP1yqxnNoZAr7gdH0FNdr/av13GHT/Qtqt6
k0n/gs01ld3AlXvN+NGRjBxzhnWf/PqJys4LotHu8X65B3iGw5FTiAZNw8tgsWfo
WFijUJKL8hoEs64hSLcYEqvn5ygqH1k0XhRd+y65pgUKoNsAM1Lw1cPRz0raGJh1
iCXRW6+2SBaUdKsLh4sm6yQBPUmjUc4I2HPEsGjA9iXv6IMtJyxE+y8d5rPbH0Bk
JIGKtrm92XAyKLKiNk/8rtCQAhi1FJgc8Jt3YCPHLR+xj4uz6n1JCb5MYWsUJBlm
DKwEVwhP6j/14atFYJ1MVJghLb4UhpMMIcedC/E5aSuIiT2TnBu2YEq8qgqownMC
UvfWgKKvGNCy8ANVA3g/ZN8A4sR1urpJtxdMpRo8PmL1hNlyaCFDHPZqvP1zIQq+
HJF9vSzYOnuhCsUDBCjnnwXhFR4fY4tryNjIl18/je8yrCErNAzFkD2ICWrqeiYw
VjTqqMaRjOhUwpoIHsJhYpueJJoh83ef7idf/evhalI29vF0ETGUFPBQ1GxqeaqU
/SpavrUyUhNsd24T81oBRgXJyz6/J8kyeG/FJef4E5q2SrqmcW8xvNv7RSmAX0Oy
O+hhzI1HQrntYIpYZcNE4dzHju0rXWBtdTWh3fbEhXoCuB62jR3MUza1wTu/j/Ai
qlK8MSgmsyfoAVilVR1wPGV03zN9BhV2zt0ms/opijwFdG/rXsnoREn3hl7ul9S/
JlWWGKenkLVqNiKEswQnGLEGxRuA021peQGr+iIi/OUlnIJtQiXjoBZhp2bIqeWH
d3jRFOwUO5phdaMC8hV8pbb0Bsrq8c0tTRg9xOA3mCL3IOIjALNehRJ8JRqPAXBJ
PV8wMqmXQOlFjNWkKm90Dx5rW45O9BAct1ep8F8O56TXiGgJAiEgJwK8VLEkDgBs
aPgEbE/xNKT8bo2uWC1ib6J3hAeg/mPpMfeu+HvGuFCNAiknS7E0nAcB5fmNEpAi
N34c0nTf97IHEtFYevHH+LDVOmZZ8xcmyWMFs4c/CjVysEiUagKXFt5l+Naex4Hj
yT3cLcd/TY44S1/t0uPQ1KXdATqkLF6OGmaR6U+katgVeHlDoWSQSI9Us8w3mpAC
ZpX/wxPq2s+3Pa+cYBxOPEyiFa6V7V5odczaIOSW41dPoG54dSOZfQpWATRdM/0L
y45xRbxEgRv1K6+JocGUoVxu5oWffQo9o3sTslzaXRrCx78f5G/3bG1FOsrtZmUX
B3vg6uKxVHSwVhyqoWOIOjNUcm59S7AaIRfrH17Vxf+A2zxSO61NwsT9PzDdTIul
kz4V4rOcSxI1wMzQgw9HloAl6N726e/WnZYdla+CtNoD+C6S8noD/hS23vBT1uoj
XawgycSNA0mnPapV4qj8fp15LKjkgl49jOzD0mDHK0xpUm3hgtzUuH2GaT7wnMRJ
BlK2FW1udymOCMlUSo23QYPhqyXzZAn0bu5QOMWv8LOdtc4yjv0Z3LXC2cRiI5Rt
36t16zZdwVcJpEJ1W3saVIKLUoqO87R7zCPBpXM4Hor4lpEGlaGPbHRz65sXR7jB
Fe6YOibwNzU2yeogtlHfiMGekIfGWu+tdTRxD/Q3OG6GxsGDJg/e6dYHNG6kneWW
hpDRPpsgwvfgeelYaJ69pFiKbK4P2xRr/vLpy4zcsd/u2eY/X6AoMYPxIe3YHSY0
h6sL66f5bJmyN5r7HSOVsIWaTtEB1NXqWR8uef13GSU2nZZnDBVaiwo9JPfp4hbA
PjhWkhp8cwoiD2xKbu2AR4mklfvmSQXxgcnF20D0jG9x3RqGS5DeqdlHqnocOvDe
WMUM34cgsdpgmNv7EL0PZAvL05ArcN3dQDdxVrT+9rKxxvoSIj3d9hnJgkJsErjJ
nuiUNCk8mDTHdM+JLRLLI/2Jyc+T7ozG9PJn3OmPN6cf48QLFc0VMT/FEoTQdlUH
tvkjlg+htvTXMneOEBsqzIit7tFpECpbpTXbQD6cBIVqGxxZT9x6XhOUGI7ZiQkg
yS2cHtVW9Xc5GSQMKdc/Zlwa5wqbt64NmmKJjVccDljOQVZvfQQcNtgNXPKJKhkJ
+UhiPHkyb8b2QxnYUPi7GqkTAdhoP/9YnX1ii3lZ6q8cuxxyHd3zEYVPniSEKLhC
DG2AbQiEh8f5DMwZvCMel1lGQEsDYNM21Ho7MpEiAQ1H4ggjnD61QLNO3g4J24rE
LhDBK61N+wONJKLc4uODD/oP/fCXwxyYDyEckof9HXtKVBg+pUfGo10xDdEYG+pV
iLiQEaSG169s0/uZBF17YAMQZLetuKdWjAly14iOmeNzRTdMTnhgNcc1QJNGmbL+
AAxaImv+Fx70nlGZxdv7G+LkwBN/9kah41Oy6jrR6dJj2YBcmdqpYHHwEA4NiNPV
rLzUfaxmGT75GS7ZwjrV2ISpAslENcKWueeicgZfXFPLAxHMt84mBGByBuSTyupy
ek9fkS7Qu9YrU1cWKgYn2P6wr+WAWAkaHrcAXiIg3HMlxcZV4iKguulOEQMmOf53
i8MfQiJgqKdiuKmN70u5gUMXeLavG1gOcmjY4Wan+Eqdp6h1oxNmLdpnuXhDQKLz
q1vE5eshhj1q6HZHMimGSZGKP2XkBylpGyCC7YfrW7gRvfIbvJZnvYmACQzi9HGV
0Xfr+0g0+McPZ1NreI+jdhsQi1aLp7AXK9Wm9my38xviuYRRl4yPRUxjxotooTiX
CTenAG5qAGd1W3qhjGQgBR0eLGR8DzkVd4PDlS3ur8KlfU/z40MDu9mWjxgpakNZ
O+4kq1qLxuNV48z3QGcFGlCAx2zxVTeYoUdR+SBfPViQfRoSETLtXmPFXOsx58yZ
aDU+7t990DnBqhx/Nr9G52xOm3TAb7z1Ckn70I9C3G6kQ7zZFXWXtArL+paPdg5t
wiiqrTSs4jJqxS7VpIf5IkiwZvO7LgNs6HoRIH/rsyc2qBvNtNg5+6ffT31kiSId
BuqQnEfjWi0yXoZ61SdyuW8xAOQGLWj4mXdzPDuqUe+a+bP8wjH31g2C4A6LS5Ny
1wFRCWdXHUJxuYn18Qh+Y2J4kD42PtVzAdt6CqieHFwqGOeHmZ2sUi4+6c2D46zL
mRS8JKKe0J5ItsMZRRIjYmjwLTL2uflkZ0OmALOQPhtg5AQBvKFJVPRlxs4kVtO7
tfG4uHjNDi108EHYNl4gZjMe4BGKWuCYxrSGV1kMSCpoHkJphY8JsBDZvAiAQ9XX
MEVvGcMBlf2amqeNwSamPpr11XR5VeESus7/9/R7i75gaKpn3huENqON1Jb/WyxQ
a6rCkkNDSVQM90m4qPyCzkjC3Mm26xjZMhoF1Dwv6qUXP8mWpg4+qXVBa9ReUjku
xK3s3xUe5gNzcfiNeEr5QKSYlb8QYYF8wcF3IGldCuKHbcJixUioQM31YfYsQP4/
USXNYwUDRMaw6KGGGPNPocTyBpgCLiSP+Qd+AiMTiV7xPIHEi3zVm65i3w/WQgSY
f5vyOADs+cG237I/wub5RGAYztZxOgzmwzTDdAtZJvUBhMp82Q0q2387FirmWs+I
y19diNuzX8TNQmt03YARQuaZi8jmiA5TkaWaQlrT91ylXUk3iyaYGnXKwQovqQjM
ke5QwbTmoXsmFErcP6vygfaoKUtbcIvs9vnxG9W+WDNh7fi+oxgABNpwAnCC7FA4
h2TRiNaKKBgzzqDPpqcH2QHdb1vbJlM3dYhVEz17yxmT/Ym9pF1CKRgnEtHZAKay
sDLbbqPWP04PqJvrCWIcsmnfJR2op0d2y32D/Z/fnuxT8kZNDAuOQLAVrlG9S+0h
PjBmGHXOfpFysiLj4TFEUDeOAHqEeHytRqOsz5Rp+Cp63y/I73D5VVb8NRdxwv4U
5ZFoiwEz3r7n+/+tfF2+seHpSX2ZWNaS/HjezGQ7p92SIzvDiItO+wKMSULbz9Tn
dGch+gKHIvwsd8qlmW0MeaGKOMcHWYWF16SYbjL9v1y9RPHI0HO9HG56DyUXVjhB
h3NCSBmB7qJWXGqzNdFTVc58081fpCUEsDCJYGAhVGX7X6Qt5cncAyGvjX8uVTMs
bXpr/AU+pcMRJe1Ol8LGvvQTqtV6bTjy94c4YaYT/XqwU9TvKHTaCQVSx4u/fP3I
+T/f0nme7g/oyE2sRs36LAS8ZmYDf/BGfxTKTZW23d1S+aITcnURA0y5o9j9lq/j
uo9jpdEemUzMnnmEilyHZavK6hm5QQM8f8hca6Rvcuvev8wqbiW2CejFcUJlWeaa
/N99kuboeDkFjGLWVDK97vR2+fpR7QahYFl4Ssi7TGB3h/RBwdGF0P8uDno+gvXx
Q0m9DU34U7ZunTCR+tlUvP7LdeaBM5uHeQVDDLRdv7fx8SaAuIGISBmPNwAZ1Q0f
sltCjFqs4zvYphAeHoTdBJYBsperu7HY3FwOYWiUVG9THMXLwK636Yb8PJDFQHZy
EwXEIjOaAqaAte8v3+tICrJHGKQ7lPWD/S53p/20ESCgQLWxKWuQfdfuWGAr9UvV
1thgJGgMSAxnUmoo85EHFMnYLH24kuTqxvRxSlPZ+YnkmKlqfzhddMHTWpfMx8bA
I3qIHLNMmroa3Ik0rMaJuLfhCgAbMzwuJF4xtAfkHbntkc+v8Y+fZZFngGAK7YZQ
q4nUe6cabFVasEyEEtXbBfYFG3tCcHv7lxNiTDun+ABz3dLXSIhYwKRi9GRttsu4
gI9JYkT9MPTxpztddJWj5iWNZp1zgRKfIPSmvoSpysMBEOSrd/cuMr8abCXXuQtn
2darjBztDfhqg6bz0lQlvKM94zFUBq94N25Xmhjh+Wv0sNFrTgiDjKcDgJzFPccE
HKZo0F0dtl0C9q7zeHabR4on/zi+oAmuVzfxcGKZO20Ogupyq9AnEg0iWxTc05Bp
37vYHhnnKJKkdFhvMVgP9eHgLCKHCBO8fEBifTlagtFBfLYL5yG1+zUlXOW8YsmY
esSTJCQ97PFfT1wXUX78F9kjKBs8iDjWlRXYWHwYB6s2lNiT6jSFzWEnXEPQfVRy
3cPMdnhGRpNrkSl4vjiqwyMm/GLM3niDe8oNxy7qb53q5wOh8eiFvvVeZL1k5tLD
HtM+j3+eCm+fhtBxMLgKqQ4bmX/Ynnz0zKM/ny4n5K54Ex39Kmn7MS1byruJ0Q5n
znuwMG4XeIMZelNIo41MCvQ2lmYVMZEB+4qwqA0jCPLvKJ3ZFZr9RM232eF5N9f3
gNUQa1IF/aVMVn0RG/Qe8CF9bvlteIvB5ai8XZI7w3QW3doKU7Gy0S7p/+0tVtgv
69x1clpnMgFzhXuqvTdMTQU4Y7aTxHYZB7f0+OkEJ0BlpIlopD8qWEAU0vxNc4pw
AIo4LaX+5wUvG3+p7G5XFsAZGBoq1MTATuN2rfEb7xmlFZjI787GAz+XDsxDYd2o
7LEskA/uLgFIA8O/6JqePO4Q7Se+ty5ZCWiWPNmeLEAvImDvLVK3xtm7bpgwx0PA
y/gUePNg48TocV43HApIJOJcoCIxyQDcwnAkn4pR9Jwsukqvim7V20aoMhqGR9RB
NW4umnrxnAFFkjRJZMMx9BoDf9sOKgm/sQx5PukCF1NSwXMIy4TXqNdRSUIHK0TO
9pJTZaxrZjkzGwk2r1xBrz9uAKiIYSt1DXQyS8ojCLKuKE3L0RlV6zKN81ckYkDE
r1wt4srYLCDVea/Mz4neuDJjbMgDjkM3LeXOQFkXOFuEgMNO21t2b6tCGkCf7Hhq
zuFYK4IP2CVuK2tYxVI3cIhZtz3cpZyuOFWQSe/MKYd/ncPYoCEcY8R2zS/LaEqE
3O3x9XmkkHckRe/8FUwUtJeA/4NRrhggjAjw+u4pV+y6w0ro1+yUrHw6oNn7D3qP
abdwSSj0Rdy3GGc5Nj/qWy8Z/VhlmzRAy0RGxwGQI3qwSUU3ezofk7B9B225oxc7
O1PcWhhg0IONyYJvDSBSdtnG1FAEy+ZNw0904Kj5lwuSer4YQ9DT7zQcTjuG2s7d
oIp2mBhmpFZiibXSAyH2Xalbxl6t2CSPHKigQOD6iZuY7Gd1h3efQ5iMaYouxuD6
Z5Y6cSJbX8iFzsJKpJe8C08vq+WVJ9aHcNKuIpIaF9Qn3bHOiMf1Ucdehmr2Vlsv
wAFlFK3ZhD4JDx64Eeh52mSpF4Ww16WQfOagVPpMheT7C4NG99inlpvHyqto6NU6
nIzZ7UClwHrQkTHqdviLoUafbYAOLpZHDtf8u1C8GHZQNIAtTkLXaPYHohJnPNoi
bOTfa+y7zNCoW6msIgPsqnDSFMxaw1l4TSXpo08p86U1OzlLBdkFLKihHs3HJntO
bfPfOkUpkuor4yWTtT6e2SUlbQ1zlkTAbNPJxvWVSFtwSVESdGXZOogbOIz8r1xJ
o87+lSl8JjBUSR+kitInNrAUWY4k+UIedoMfCF2PYkBADZvrsQ1bIchNmwHcPWkF
FHXvCeeBkmArmkcHq6DIbxGjbUuXljKT7YFCNbdDleYtCnQXHv12U+cKhqgWYEUu
CzebPJc71XdH5DKxB6YTBcLDO6IwLyu8mZl4qFIQxgdEOGhvIaoC6fCfL1LutXS2
1Sd1hJLinOoZb6K3tj6TiA4KU9wUoW5NPHAoKyM46zUkoas6cQJECQmiJ6UpVHzW
MKP3YjyBTJJXVnKXdvmKow1h6DD6VoM2LFKZzEI3OHz606CtiByHS8/QnczcnYwC
ZvLTmctxw+yrY3gAkLYlEEYloit4w5atz4MKAer88g0Jkx6WOdkHRkyeQIlMr1Fe
YgxrYi3hdFcj4uFWy+hYB7J/sNxTOKQ4xMICVqwQNu7ZDvWWOitaY5pyDMLNzY79
k0RAQnutlcmByTZlv+jQHO3EMjnkpJQG/mxSpjlAjDTVf0VZVJXjDtXD0oDGlLpZ
2gfvFcNB/xMhD4JZx7CaSQu8dmksy6tdy0sZLTqX2+0tnlpVHyhsoVxlTUzVp9zW
zx+VQULZUpuWDREkF9KSndv1qIIG1p2q6g1hQ5KejTN/h2xg0VVZMFTkBCPVq1XY
mleP4i7ToUK58lEhcEjOo1p7rDY3fvTb8WV/nbjER77vIHI6d/OCPouxg5zQJOuH
Yy5iS51KUbxdItGJDE4eRNlOk4hIIbdzZGgfAch4P1bTkxMz9bFZuiVxO8GYTwwR
KVE9UeTwEmj6ZMB4YVYk8Q60TzN41FZprQIqCp20odUik287sLGQioqH+by//TGi
HPosiz76ColykrFfx3kVqgwzIFICeeMHt6uDQga+zl9hrYEKYjpVCxVVm6V6RdfT
m6PCBHoU2cfNnwZcEB20dOSN2EH2K4gYjPiaGa0y/VQCSQVlroMTE6mRK2c2Qo5E
tFVvVsxYiZ7e5wKy06VdOvuePjCiyaaGfuKDDmEqEPSiAY6F4LpEWA/9aecf4GA7
ehqxOIeoWDlf7Jf5wgerAEzG83B2mIrMqCEj6ezdQa3AZXMpCA8BTsI8s+IqIGG3
14nvJB2lo7UOvPqSwrkNQnyXD4eePXKkp5FINi1Fu17F1HqxguUyrJyiCvXzntY/
TuRD4qvnqPjX8d3VYhpw78Y1eEwud4LknRgZzK8DmEyWzVz1nFJM8G3z2eUbGlT4
Ia5MhHafey+IWmrK834xN2UcDCfOTM+gDAsVU9TRbCEhrFMYjqMqzuKZMDDeA2+U
w9O0C+bky5AZwAx5fYg5jz6uDn8BebV3CnzjxxtGIGxkFCnWvyffukMO0KgUzUOU
Z30JhKdTERdE9qr/GCcnnB5c5xthgSS5w+sCxW7svJIRTB1k8F+bROt3vMRVfyIf
2GAKugwkestsMsdDat8L4g+hyowN8InPd8eVjJy+9eDmn5bh3oGP2T+3+rLjJuZX
Psh+lV6x36HBe+39pS/eaVApDuaNybGXcM2FFxKdVgmSM5BZu9F0TqwgsC8Gioeb
c7saYAulJyhOoj2FAdFrpiVQnaT/iU39Nf7JpwN9u/zXRA3e6K+OAbKmpWn1b1jW
rmHS3jLjDXk1uE7VoZs87O27+2ola8c4ejbj2IoW7/NrgaPuHD+rFhSjj+kRNIRr
CvrDvVwHvhwn+QzsaRcZRXJaqv2PHMvP4jfD9/REuahEqBDn8nNSRK0ftdpL673l
tpuQKrA5toLNSixOkDtp9XbPaVCex0F/58lH+0aCO31tSMv9dVoNmLR9rAnik40u
02Jm9wK5l+PuEAH0aHjGw8jaqMCn+FQw3+Gk8bU7L0Aq/e2+t3ViTA3bNcHULMK0
ZQojtyKH4G0HwsRWhoDb2mKBOfpPFg6RwZzqLZPv93dzZWQdVk7Glxu6Yk7TZzll
0vk8cUzH/1EwX3jERIOOwHLuBs0rovXHlIU+KVMg2WByjUtyjOJoXMtG7B4ZKqqP
s3Gom7bA0wWiTsU7m8FApPnqOIkNc+krIJAugcU9tTrgdZxhOncL03Gl+W05D7c8
dDzrGOZFN6KfY6JH+rxJGbyDrseBXXOW4DARFspsU/hYBUVUANJSJ/MrXcDVVqOR
ms0oIjZchGeWVD0OUYyp1LmYlXY/nMKQR7AiOvIGaL74zkOPDA0dbYX97Ew0w3YI
7XE6WYwA1bk+E4m6Yx6+sPF17bjYYLctO3zpq0VcH0XFSHsGno9ICAX2AoRr1Wtr
9rlDoZ45TQn7qqA3jZKBgn/1igJsur4QYe/3CET5GaN3nAOxHxKtv9xlu0tbf2k8
K6FnJWQnPuCVTEVu2ZTD85KhETmBTu0aUROAiBZVWz0ul0k5VELtEJGkCfyZaCRC
2h/r/14TqT3X9LtQcMWDuBAflJBLFES/sPU5qVHu9fDmoNT87JsgkYWXRlMHR/fe
RjbHtJnSyqLcqJuYNgll3d0EOcywCqyUVVJ60CnmJLpAXnCy2VRyzHVF/s0oHdsf
dSGkAs3Bg9aYy9KBhZnO7iFUZxPzAD2yVtenIGZFXkyP6TvVKny5YaqUHhRQRst2
v9e86qrabtA0NJ8mvkv2LwHW4skoSpS4TFEV1rbWa0zOcvBz5TYpphvCYUSpwHWG
Vl51AVh1lN4IfG1ewj93A+H6/HTuagDsj7h+DpWJ6ggM2FKZJr6KS/4hqbM1/bzN
Wh/ztLYXdy+ktdcIz0exT7iJTsjS3tgXJyXvG4NqpdN+cZ51SMEsgFN/VI7KFlpW
3R8oA2aQKpxRdDR/0CIiPoqRfBJgGVL2xiPaT3/BF3Bfj3/Yw7B2GFWg+iCNbQ/N
JdMsCZHQMAKEoRL3vSlf+s+w5/W6zQrAJtVjoztAHiQygLu/jzb5pljtyLTEGSA0
ZrqdpVEbMLG7YyBzQmp+xGQHiVjhDj4KLWFq4GvS/5FWaImf9v5Sjuo1LtmdxsoR
y5HYLq6y4gIy9eWE05yO11WTdXOGnGsJeCsUDe62Ph1LtaqZUHAurUizeHO0sUa4
f3dWAqokbaAxYoyhmZzgloNYdo97hUIO+z6Z0HTb/lB8M6T0y7viHr1mtMjnPW/v
FhH1RWUTo7fd+VKgZ9Ja2zsSosJMS0jKKHBVZVKJl/Tx8g2zP5YTjwRzbi91eSBf
bkGQwBnJmcQYQT0igN/4XO6oO/KcsUwQSAUFpM/wzrK4uDB/FdG27zivd+sOJTFs
MoJKL5+pnLdE5IynaVrgCzV+QT/QphQHOLoUHUA7FLyMl/zhS3MtEruB3cEjyGzH
F8ZK0UXM9c4waQ6JnoWPe5uxuttskOdZTfVz6KqYFAaYS+GiDMUp+B8TFDYHCzUd
IP16haVTuaoK2prYHKiiRWUDzmYmNvtkRXhTA/GTGK+ar1l8BNYLVYPV8Z0FcGf2
DRIyKlx0SZBg/34W2v++hzNwhBvEieGrHNOJbQpv55apszIUOZolcAXaW7KSKkAg
62N2crBH7qBjtpkvmG/oK8vXRfW50fwiO4iXdovlFHAxWgQMCNDOgwOzZb8rpAn5
5z5pP1657qrjHEzx6ID81JKSvIZjOOnL6CYBX/QNsbVdpid++ej0fpsIR6u+pGBm
PQnjtvUc2/Rq1oSENu6tK5d1ThQkQ7nqu+AawLZSJOOwUvEe0ZJ7qmzvGdSQLagy
nFL7ILd7btsJvDVo87UJXOk0sKZSRFwGiomIqEMnrB3/LEtFH3BIkdaPzblcl/AD
/+UraDm1Y0tSNJuarlQB19bKX6mCtTvrOtZLENaBcSUQiOkMBnC/DKwfXi91KRtE
wEpAj4gViVwMJXPrMiymSwMA6qqW05090rjgQv7/DMs8uztVPJHd7yN14tmU1/Rd
DO7D7yEwkHuVtmPXfKnWqjRTMa0dHk1QjWUe2/dqdUYCBQJYzxZ9dkv+4UyD4OUw
SVEpT9EKtB9Fs1rkiAgTWCQYhdbovUqNln733twRUPKZ+WSAq/vLb/wB3xF+5fGf
ZVS/qSoH2Pfxt7h+1G+wk+niUsZizIWtn9yjH+JEkVRdb77ZHTj+EnT2WdX4OfJc
qI0NwC0sLVUyz2bQMYuq4e9Jg0NCTfObyTUqoqJJTovSoGQY5xeUdFglfsIhE4o3
n1+1O+3ClErkcnQutmge7M8TL7GvWwv4/eUf53XCi8S/eRjEBuJMlxX6/MKBp3ut
f05vgYilw5gooyyWy/n7V6foJws5dahzZA0ICDBXZ2H/njkUuJk5ihJqPVYTASLf
yzP8jMG4T25CYlDDZVODm90nUg+0WCQ5DXMzgNHyxHTtR0d2YMHdhXVN7FW0+hHw
sW4NSWuWbROHUTJ1hBHaHTWqoGluEusxmrFiXaRSUzgp5d3TazJYj2EnbS6zJ54s
uNcJ2DSAxheZtft6cXodb9ckwntcULKCCAgzAmCyPmIyXY31t5OI6SDmh0lXMnMG
WnHsd/GVV9YKWpX4oaHhID31KRvoYBT+s9yyRXZp6Uz2kdgjAjH0nkNoIsYKAnIh
fOTxcXvlLf7V36IQahQj3utRtw/Zl0TsGs3bfa/ukgfLgZDl7xgZMB6tVv10qOXL
QiwToyVxmE6y1mA/w0tsZNWwe3rYOZ95Q9wybu7tzHAM58wNQP6CWuO/PviNRuXI
mmZFrMyvV9Lq//DjoW7mPoGUx2nWO31F2Wt8/gUlXW/SXUAN2XWIICnCONWGXfG7
scCxOgVphXXQ3G+2VhzZ/QiMvdjDCj2OcLro/h1+eSM2CsEXbvlZOIPZDOKUh3t2
Xw+KmJTPcaF7hhxAldTX57QTDPy1gm9sJsGpjRNppQbtUxD8wySzfRduULAlNmb2
y7zDacTJ2c6HPKAV6iNFwiq+O94oQFvk5f4MTDffRZrtmqm7AWjw31lB6Ny0gVt1
FwGT07QmNGfY8PWUjm8+yGze9hFz7/e/j6fj/I3A9SoG+JGCjAgXlnLdvu3Qmws4
DwbqNL2a1JesvEQzetQY2l3I7KVdsk3GCIntl6yEyYKae5U2Nc1wlS56uOPrB2cL
r8UwtDUrKddjQG4O+Uj1qTOkgjnPGJSiGJAzQG5aUtf1thOigoY9Vmed4zw1rCgr
78Y9VyBTuVPAAOIwGgds48en1Ck2plZu2lWCR5y3M8wrS05zhHG4VXV6Xq9oNfNv
e0FB5NqGWD5TFpOtay9CYSoW0S5JFFkIM4KhtWk3YlZrUEw8miMNje5rsqiP0hLb
Zlp3OrgZxKSGPlrRsuu8AhlomaIRS01dJBLQyIAXEO1vu+zmhIqPlcf4p0oT9kDl
KVAbzo1oN3zK903DfO6qtp8XbIj5crARhdoFydvlVytQP1Y5EYf3Y5KXKG40cYFZ
tWaWedLGAXHrbAMRTQUFIkClRDDN5vPtD9FRSiTQ8ElS9q6X/RCcveiw8DT/m9B1
jrQNS6owuB9isDjwpuhaEvVrwOuRkZvrnLAXMBMHa3fu7bUK15neFCEGjv/glq46
B5yfkXn7oHM3L5UJAK8/vmWs5rrxM7j1dotVbbzr5POMn45rJX4SIAAjNkOnMOhB
aPlPfbsubifW+nL/yLSKBqXddDzj5TiYvugWRnrkFpVkDlR87TZ/HCWzXvdaq3qg
vGNiJl+xEGvbxQ2eyDa903KTIJoEZSdgBAX0cqz34tdKZ14KBu5Sgp/d0X3AO3mW
Q2ApkiTIkvxQ4QmbWQQ0QBMonsNlM9xZ6z8XomlAeQVQdYEWPlTSRkY0eE6r2Z6l
gSbxSO7zksumVNBbmwKATxNRDBNVySq3y1hshR4BiEig+jLooljtoqWz6YMG2LYM
IDv8jkGDDI0Dxa7sGhYaumpjD4kkv5PMvQPHXTrVT3wr7VEGpa8D33aJTFmyHNS4
t8JZGo3hiqKby45tD8wfD39OGosx7bYFsWUyxqdd9yqftwWRZ5oKpKEHf81B65q6
WBrufa/+y2iobLYGY85dfWj8uln17zrP3SNe+ValEV/GOprV5H+BxVaZaWzCkk+T
I+61Quz7h4NsM1tNJQmDIhIkqtGoqabrMB9paqz7O6uBnx5h6yv8/z7/JPaTGN2I
2RejaXYHVvRMtcp0LYpzFTyw/PT74PE3knHr1sB40fJdwCWA/SEQqWfKmuJTDQ4n
5dM2wN3R81RZgODuNA3iGqjWE11Wd2bstatm0JR63+cRXBus+Ja9OwkeBFG/jqE9
goBlYHjYycm0A/+oTx7P9Kc3hRcj9tNvs9J5enndxz4wXXFTEP8PZNWNXotf3lDW
2VgVYaymlnJavoqNbTiOGQEwtwM3Bt7xcZCgORYXACSNKOazOY6HgLG1NNNgzWx5
XZm0Yb8qA6F+Uc78RO7xyCuBN9nawfqI0Dmg8rzT5dhiDZmeUoGdoCbsggj367hb
5D9BBi0N15N4qi19ZkdrryOwgIn7BSSkk+bep2s/jDaAAfnR8928UvLtusIGpT40
GD6a8bRCNGFobzI/1PMcopQ9IOgGuSbsgPyc/XQvYsxVE4AOGs64ekCyNOyJiWZo
Kv/Fae65vv4JVbNnaH4I2zGi1aKk9pQyX3bKvS9Ao+msS/OyTByOcVZZL9272p1c
mleTPloDu3qKexy06vb2i5E97vsRCXRthuQ3i5ZwO+T8u6Yo3TBDfvr8aPozvN56
obdKASmAkL2TDfkK4OdeM4HsaG38A8aEEF/rDw3YrGHXWtK4DKGjnbh4TcP3eNLm
xh1fQeIcrY4QJCSMbwMfNDp5KEC977Ls9rcP9x9k9NqVN8d3eshexxDXUcayOOco
BcYTVYvglCQlmmAkstO/2km1GcHtomu67AjLf03lVaGKg4YghKCVjV6cMMW2wx1S
diRtpTtP3j2fYjwC7gt62nAPWePeO1Izs71b14bN9di6PjFP9uIpzbkyp4hZoyvG
D2e4q5Nesdr6o9yVY+Uyo9zgaXsPbQ2NhCX/t2Xs3kTHoWDLT1Bi6Q3p1ytswzBz
hdGJT9DOJXeH2AlwRb3uXBw8DiUC2YZqBXhQM47aTyvFIne2fbgjZi7xIkKe9FWD
LBhAWmJ8sN98N0K29TUVqPi0jOK7JISBGSGjj9AZMuOw24ZabArX9mAZI3byoI50
HUQCjFrtaJuWWLbQy2MG2zQbJeadyppwAPFVuPTz2GfKPyikO06DNlrFJ3DuMgAT
9NLkFykEondlf0lk7i6DfvDi4b7kNHt5HA/CntOl0DhoLBydOhdV0wKx65N9VNxb
V5k8UDHJrDQ6DmTJESjrP8c9vax92B85yOhZ1u6LRJrUrf1r5oymbg53Tc491w50
tJUs54/sJv9/B+6JM9K4wrdNqi3eGE9qWskoVmxUpR4GMcVpthlYhUh/U74Oxblu
fXOUlu0dXzJzne1VF70XGu/x9dcRxAkRjYFHmoZst6FPpS6g2tqLlyaXhqAEppls
S6qC7rKb80z+ohgA7jW1kyw/wsxP4vTpPxhTXEs3lJUdlypd2aa7qdDztEX/Cilj
ArsXUETzQrs3hHfEh5kVOuz9SOyqqrFOpq4C8zBEEYIajf8DR5YapktAMnzLawa9
Nkepi1J4Utm9VkF/7R/juEYESLkj48xWosQHrzYPcT5teTeJI62pcrd4EzOvmZmn
6IcjQ03kHu4v+d0re9PJG2IqLENbtGZoOR6xcnxKNxzm2GhURwYiyOKAXrNXmz6R
yVNjj/o9k7OAYTDkf5T+xuBc4nBP4k5sJZ3tP7dHfnw9Ulh7OsJ7paRcS8FicVcQ
7a8D/3Cy+trDk95fPn7EpUqFPBN3qWn9tWgPQrLSL8qTrUSOWFvyxBl1QRlOgSVX
obRcYr5ANtJOoIVXKX9veJOjUPbfKMoJ+eKij1IM99GK8MLWnkrtm+yTh6FFtgNq
VNMEozvtxN4lp3SkKcoFwVU92MkR9tD6xk16C+xdKqh1VZX3ur9tbxKW4ZIE30XY
0SF10vvhAxOTz2yc61w31TJ3DMvTJRntiB8RUkV1OI5mtl4CJaMDN9dL7i90Vk/h
xyyTLpUjjKkxcEpl1/kRIE7o+F/Y86Lv+dOxxt91K5wxnwCnwE+f1GLxg3ncSpWf
daCebfzMnCCm0sCgqfp18qpd8vxJ/9xvPxM/L7cWDnOGaeo3tX8ITKHaEEk6u7a/
H78q2fJw/vDI615cwOGJARQ4s5AXVG3yHfvEVJQAZ3P1DionpoDEuYwyNmghfUh/
EhA7X5+ti7QZ2+MKDRhAOQwj32bk4oKA39duvayMzs+A56rTKQ9REMkyku28eMkW
uVAc5lV06UNnZ0OQYajah2zQjydJqS8/NDbSVzgmbADPI4JZwxdNp+sPUBJijGGO
y6QKvASfC/9P0tQ/CJDSPJfTEtiDF90kiq38jl2QaMM/ppx0kyIJKSy8NgSQ3jhI
dzQnP3s9fNUO4SOS2UMxVJ85xinzbBIiYEkkTHPtMXm/Zx+mjn0gCtIi8opdyEDx
sx9GD0Ho6dF7T5qcA2l8lOC5jXVIakCr2qiloztz3SEzh/g4t7Rs8J4M4WPoztHS
WHTDFlxV9i7XEQZGgi9rtGVRrNK66GWgt62cw5ZFIIjC3e/JmzQomrjoYYnx6xHZ
V3SQNL8g6sTJh2GHAlDkAnOPt7NE4XCXWsUDkkbPhtMU/u23Tk9B1f3XaACjKly/
q31AeqDXk48LgAsFghcmJZdnOtRP95D/6mUJZsg7N++B786RwpNWgXK+XkSBRyIJ
x4fIBphqlk4aTXR+rOgsbhxUNNriBwHos76QFI85+pRx9x24je3wq7TTx2R1yi8L
KnH+Dxa+VC2VpdzoLuXyXZwD28P0904H0AE8IpblfDcgFATti1OeQ+eF6zvb+s3P
msRA1FS0b90QQZkGLoc2sdH6Xs1P1Rv2RioTNbU5OJmc8W/8STop5bpKZTRq2gOx
e2I9g80GJcGAazi19V+oq6M02+gisN+Rj7oJ6Egk6z4l+GmA1rsQaOwQIhdqxGTd
AYD0TckxRmvpOCEYgi25sXmkuvqn14olQqRRUyBFginrwLXCxQ61xi4CX/oLZh5e
ypckNrY3nVJmmKfFVZoqU0j77K/oopUoVbUtiwg6H1pchyE7N0lnFn83Wq/TQhKE
KzDWkDocGJjsEDieEOYW9qOgyixp80RuIkApnmVOZMHInx0nQx+LRH/QiDTFV9xD
jvYpfCdD09PaDp4Kyq4x8krvSuUBxyNKy/xo9jnh7C7SOkMoRA/xeuTmFqGc5QZQ
3K/7FTD+8CCvJKq10MS5Rhq50IZRv0Pasbs33Jq7gwJMkzOqR9OGDr+o3MF0VmUf
Q4gR+esIycLkjKWkT/q4/PEBjgsNdmDQ5ZTBdJR3Oz+uvcFmyKgL3NZBH8OJp8Jm
/C/vXTyLnVDsQd9oUyU2H/1FEG1JDjBY3mkeyuVDyUKeO4ZSm+JMrbVDcVRpCs4/
yUZfht4D3iNpGaAWHbI26ItNHYJaXk+iRSACWFtS6n73tRcIAXSsW/uADa+mAhen
QkgE/KgzmyldXANpxOZpE165wqzMNTXRTCMCdfQnP0KuG6A4Sf4hmV2dw3izPY0T
u929qyd7oZ7yxm8UdAhVuX5r9OhFBE+pwaTIRcojhYFCFD1mdc3n3RHNDBDiKttI
1XTSqLTkmYgL+QcxpSikcR8CmijEp35i8vDg5qMq0CuJaaKvpHqDH3qym4m0Thuv
coIvy4dROvwQt+58HD7IN0FpPBjAb6OqMH/WLnkeCXYOhjRcIBf1CHQEB483I7RJ
UQy5OONjii93GQXmSJHnmAtdmxP5SxlGjTZ4bRFjDDwM6o0B7GVp6qNxvRRcjTAB
LSPLs2pu1EOqhnSgw3ZSeaDMHyyED+o5Oo8XMzHHYm3F8JOl5M86Gcb10qqhnQCg
w0ebBsPXNxPy1mbJUaFFTBMRxW0MXsRrE9DMktMkFhHHUmxN2k8axzDbKHD+8tyd
u0NYU7Nur+hMWnpIigLXB7iMrMjtOkjbKhvG97Y27nm23bvMvAMu24K+qVPwSfRo
YFGf54o4A+f3A4WNI8RYJyeeyLn9MqzVawDWuy6rbVMFaaYkR0Tpz/5s6wsmf8A2
R0rH7/U0tIhdT5BfJMakhh+CYRhuRdM/v906lg60TVFrzW3fNJinP4s32Uh25gAM
Qlbami9uQ9ouRGsfbVR26C+JKdUVyg0l+TA+B07minPScea+PPtuYmTg/SPC9JEM
rKtGqM5F0xAwg3cGkObZYLjdryVDuesnv7DEpjQMUo9HCjKTJOUPsywOgACzBBST
C11g4IvpO2b7+n+4Gp6efXx2AwB0WbW3+KMVeoGBRbHwP7tz4eJwWOrYDS6zvz9f
d6d2hJHkjf+QedoGRqdmrUAzu2ntUvApzCVIXKHIe4EIQWl8FBZ1E5+fo0pqbJ7t
RVjr2qcQ7sRJp/c/KtVpSIzz3LrbEGtzv4bKQGBBqisFz07i+9YsKpuHS7Zg75Xz
ZExG6wWMZuuKZk1ggH1lHq34uA2530TH3WJBbdpB72ieLlEYkpmPwbEUxtnzYyP/
Zymk4CnuUlNDl3m9pqX0iAxwkkKZcpAWp2u9pxw2IwF4a8B+gJnvlqwyjj3/mwrP
FAJEe8E3yLCWPJ7b7Br21DNYUkQNUV2AzGnlkRo9hz/IRtilpj8KbyBkFIuZCmvB
7CFbt+DThw+oGj1XoEWrZ0tyO5pfYEQu7ytPRQKlESmS02zj0Fd52C+09YNcZR1m
zUeVZmIVodxNpfwv6CwuQlPXUi/7vovjTUhAx9SLhpbae5n9pQPTlj/tmtu2Hq4B
IysDJzawUoablgHNryDsLzyp747jUOVnjbZJ0zNbL2WJdT9J3tTN1ZT5XRsRQOSi
O7VTG6BEzqMnAdnjQ/FCaU67AAchgLGZ4Il0XaGmrLuQ5MZZK4Puza66PXwzcOAw
LxoZeO0sqLZRzUVCFO8t9b9RQYRYCIUDJQtWn0EIgN4on4aWJAeNYIioXRIOcD2O
EdudNRpGor6O7Um5K/8YmkBp5pIeCeXw9gYUoXc1icKFVN9sagcRwVYusi0w/2XX
3WT99pYPrPF1eDFLCB7DbKWHyPtRS2b+RTZZyJknlh2x2t+m8Ua72NQv1S+BgSxD
+IAsazycql/x00NboM80Sk6svbGeDKMw4UP4lhltWoSEMFt4bK+rI5bfdtSoNVF8
0ui39m+uYGU6JX6UcvbpHr8JebCLz27AodFFqtP5yJMTgEi6eIpC8bvOZyI2+hqq
Ch6KRXOJ+r6Uu7rNskfdcn5Xn5RPIyfmZDWJvymVLR/cFKTp4jJ2ElP1+Ez0vkT/
Waf0T9Z4Bvwrp9CI0LHFpDblQoaX2MWUzLaQePtB1sHMi2azwYRvGVezt3gGMAzp
OHd7Fh23qbwFChEjbqYQh86paIzFcOX6/n/bVbYbiGQwfcxnS+RIW33ONMQvplhs
9u4licpuppeCO00OhEDWsASiwGbF1T/VbYiCj7cvHiJ5cH56BUKRkq+lIy/dqOXy
icmXmqLZq0G4+FuK2iai1fJ/a7/hzQKVHysGs4EX3rniIJVEYKSCJOQFweMTZzA8
oRPQidemcTphKCmfbobGfJzJl0fdEt8TdXT9R4VHME7kVbA2Q7a5aGB5Hf2NYoGX
3KZ6KWkIIf20qZPF+QXa19OuFovu57nber62VZFEY80aI7aEw0cyjAhrvREmq1pq
OS0Gmj8LRPdRsE3sk1Ro9WNal4b4jc+udxOKCFfyPW2O4Bmj8pYsJUvouPF/uxsN
14ewOt8yYYaEz4+nZMeMtdz3MAWINfluHPZOCjN1bqOagYLBn4OSc7ip64MC87m+
CFTRqFQWj42b5HRIM8HGOvjd65G5aLS91I9/l3u7UtzWvfY3sapFoENdDTLHvTpS
i0BsDRuLaWt1sORnRADwILXDslp91FxpdHraOrd7Ql0Y1LvjuMRbb6H5SA5Awkk9
Z7onHdbrkyJs1xX7pBLbD0ycbXBhCDlPPDI0U+xfEIh6THiWCvCFBglxmBlZNRAU
HmtEHu5c/eHrhxvm6TE1Nh7awckTOeVlnD4jHS2YYVPYbXH9Ux2vNvgYFeC+yxOo
UOi902m4wlDtkMEUB/tfpPgurAq3RyJGh0jApZ4tQ1KjqAFlQtNPI3YgkJYguJRF
jVqQvQllOBgB76YJJx7gCDtq5C0GmTk6DDGc2wu/OioYPTl0hTuxTPKIZGP2Lky0
5ZygoiiBnOn0VKV3e0gjnw3gJyY1JFrfQbEYbDKDWSnUQN50FCPGQK9j+uLXCfRl
AqX2AMFK7HdM0/hiSOjD4ZZis5tQWBxrJHscPgkW7rryF2/ArO+Edg0aD4DJE+nH
/IOWFh9MW9jFmHhy6WkC0oeghk6ZxhimY2NuGz3TkHsWxnU3bJlG8W0NtZLAoa8z
qDWAQe9NBPbjr6IhikIT2PgW21JexIAlzKAXpUcJZfT2+W+50iaQl6h9R/aAnIFP
H9JhH+GQyDG+VmpDP/VTp2iYaJ6+OC4RRwLvaBD0w6Ifv+73Ncqte/XZ6y6QbvJG
i7lk8kMgIBKMzUraT6cnVralq0hDqsiLhic1sXf43wsDf1b4m40gFHl9sFGTVkRC
/N6Go4bdvgbabQ/Ek+/humTviQp47XYQMAwh/YAVvrQrVU5byckXc4ZHfzgfbG3P
wRNt04pCvpCulLrmSpbpgAU6E0N41HBJaEkHlAaXs6MUKdqT9GmA6gwccJgKk+qZ
Vlq3pGnhvclImTYJxgpumixMOglxwhjuVe9D0JvEmzxZprrA+Wxj7lacwMJWZfD+
G3HrVjK6pi46XmjR9sUred5oTXJ9yKVmE4XVOwvkU2GzoqsdKe8dKrVwBxMisdym
zYBaIH4zQdDP0LJwIiFoJZiiBoqMZ5hYIxq1DBSzFuN/MKqGbsOxU93grJyDx6uN
OGe1mv7Ei4moAFREIYClhw/sMoQSKPnEAhu5N2JIqYPfkD/C8hDUjaGpEsGFiPiU
Wc+ST1rQuhhoMfH0VCW6S2CZPmWz86f14FgourEY+HOAO89ysKEPjTzJBHT6hfPE
tIkKDWxI2wrZvnLCUlqjC+p5xh/Xw1P9noMZKv7iG+kEZCYMWGTmebzk5+5IhqRg
mD7QlBAwSuysGlabk2B0WUQKW9tU1ohYp9g65ZvvdpIfro6HHYJouNsdrByccVU3
HOjjV6QNNJExNl4KA4jQkNLxU4skHyDaJP6GhMF09Wy/VaLRcnbSekm/wpYEgEd6
K6rNOJcujd6G7JIiuOAPV3S6QLWIwvEfLBXM6BTi/Cn816Lu9kyha8mdaIreDT9K
zwVw+8QmVslGfTnnU2x2zbZnCYYRToWPM9iZ7ZdUyodjZ1KMlmN3FFBvQVcbXVlV
ujn+GGtsKzFzHKxLQPSPwSygnwqRpEYthQUFOfVqZ/EjkK/+f8XYXf6bLpBok7V/
KxwBjSDa2W2xofiVGS5ewvU5FxWUx7/udKl5GX2tYcCp7KRUAB7fOwgc2ulCAs1s
pwmo4qmn+P9mwfmnI5yCTwd9p754M6gIf+0AzxL1xTrGiXpy8VaqYAJRBT4koMbi
MCLfzJK/2QOia+XZkqBhqjqrDGUk+eIOdJbhLI8hmKVwfS3z4eNO1/aNqlBKLC1c
ZHJrKSwjAXEsAKELRW6pM+z5DTUp4Qsg/ZPYf94Y2APS4LJdNMFZxIG64tmH3sC+
CsNvebmGpfY3g3juCc7xitNYFc2DWvSFeaBfPG7oTXpkKdOMqjMBgZdZg60jl4vN
1+dCSWmlAaRQpp/TBqCeydRMoPG39jhNzzWYlpvsPMm0v5vajIy5Xgg55pkqzlRg
CcXd7iOqWhqiLSqx8ibKSGM5r5FRnJW+vOGBw8XCJJSn7wvsI3HZ1EE6Azrfkkvo
3i/iXegoLAVsBzAHqtZ1sx9jVdLKM7H7RrnKbUGankiF4DYRTruhsVGMa7oPj1Qt
jMwJffNM26P5omRYqajyqbilmwPrD2DQmkZCfdSqY02SPzrLWIcdmQIBKewOfuyj
BeaCtj4IaSlJ1Qse1gBXXhDf8lq38keoxWj6RbL+XPf4fGvejTqSOy8s4pFGFSl+
D6IzWKV9A/NCXT9CabcM2ee1T7wLIcBfyk6uFvidFRGh+I5uo60K0QqtD/JsamLp
/fo0yaUtBC1LUE7ty7ynJ2j4X9rfjXX6ZmxWms530aNsVhlkrPhweQVDcaIEa/bw
jRlzkvShfoyCsUD0TdaskARoLnHLrCVY+lteWwSgdGE8cqQ33uj0NfQvJCRjasXV
dtX+ERoYDq6HJbLkkfQBN9pM12AyGySvIaiHVHsAlq8T9eRynFUvrfmyKK1abZWZ
folog9C7IC2XeLVbKsSIWnT+5sdMYaQH5ni6LVMyvSb9WGzZqDBBiH95KYlGRypi
wlCgdb0jNfqP2BAMkkWUF0s70/jCldOwcCImEsF29DrFE5WuasKCy2DCvm8h2NR1
r7DG2xpkTtbtnF/ao7axbCmQQTVHQLGJGnWlhxPxzrSbpOOli/ZIh56vPf4PeMmc
tdyWs1y38R84+XKQ9NV/AbKfQElQi6JfMXIXeQ9EqCDXdUTeXdwV0tvPyze5PkhS
mgAh5NXOeeLaLYDRRkgi9ChR5mFe2da0D6/fuiQzqOWUBYm2iQTjCeYEGGvoH+Mw
ilPXyVUcRoZ25ayDaO0+1xb7YaovSTrO9s8QV8JnlbfDP5bTaTwOPQLLwl2casL9
Hg9tqeWKQNwxnpJPk8AxhglUFDP3fc6meSUuNwBOrLj34+CntfHnn1a9DBcfrM93
dcenXvxqYo8qsNOCqe3g37dOlB3bJRD8qTMZQleOFo544OWEr88toH00RvrdoAdg
Cjct3gu7CLK05Fh26KRTMPzd/zNQ3cEwpvn+HJT2yzbWlb97JtMRjfry230xVFPA
QtRg1xeyPMkeBq7V989n7AgzWz61Dd2P7HDl7fm0ibY/P2sdQXwoMkKvKDdJ4zqT
iwK+5cneLDg5MHiHwYunjFvoiW/BnhM01Vs2NbxuW5KS/Uq+552Foi1plcBN+Qdg
Hdrxg/bY1l5XHqSD+hU1irrjDv53LnX9j3FUmsUepko9dH/YAZoDLMPfXEY0vJOf
8MOLc9MjsPTttYbSnGD0rg9ftsX69tuvhpCwYokbTtdG502ebSZbEDAxr+2+ovgc
j6IH3Z6+PQ0Jzh+4sfnlGDi9KqnM7WaMMYGbwtnEob+WfZceiQRIYMUE6J5753IR
8r63aZrVwrj74trxH02GwcUeC+PlHPUjQeLX2upuYoxUD5L9jhQV7AhSzplJcNXY
h9E+vF+qppkSEma1MgPBc5gB46TsVTWmcw4cBtCUux6R456tNlqkizRsHKf0DaTv
ZAZUQyTQ5hcJe8IMmoQUVLrclEz6KESu32XlMbO09TktUbqjKNaZqyR6DOfJHvX4
ZhHgHofZXN/KDrtvvRjg11LhfEEi0toLkTE0cbkfA7nSGowB3Tge8a9qrs3zT3AX
hPuUBTwzIIa8N5hzNeQMWP0rqpKj3bZNTdqOcAJUnt7MQ/yqiNkDESRWDdiKEWnx
mv/x80i0nijpjb5531yVzT5Bf+E9YafEUr4pltOEcXwAy8TSMEP3mEUv6++SNyae
oo+1cnhubSYrMhzz0j05sXyp3rjI/awR73Oo+37V2fT0nWIKQ1KerFO72xCQIuDU
ULx8E2836OW4YQVeK8yBV7u/Xmgb+qDrw4W8YiR51hjkXrDj94SXpYvT1bZddH6X
JfVnoQZRum6zYjFbWGB/Qi2RAkclnF3PHZ95KQXZ5QzAcxNeonZieMjwkVnQVa/j
rnSBgQ5Fbxj5vkEQqmJncgEMLKCv9/mIQrfEcqsCpLQPb/+gKahYSqXs02l9btnZ
+Rej5k8n3PkFTEZERhYXV1WXxz53rmi2lTVd/UE/4m8FcGIIc/oAvYpZE9ZdDaKc
WlSFfKlJiT0oyD26Qondv/tHMDsPdAsPYOzamSFv315llhhn9J5UEpIIL3f0+tw4
WOOym+DAaxBy1s6SfHl+Z1tMTDkdNi/4kkPCk24vKGZx5eStzeIMRmPCc1x5Yyu+
eHtteQVs+vXSKTJZ/uQxDomOK52wmE2ZjaSpUOhvyxIYeZBYK4tIhWmTnB2CmU15
nrj8HcvrpnVsGborSKET1awdBHCQD/qKJ7rpjvZQzrb9RPMXQl5GKaliW6ZmQv8H
F/hkpIaKh/BWhSd0jjaqQtYH6fQS/ZRETKmsUZX9hd5mcLr0CsaU8KCDpCifSTCy
9BwMvVZ25sPoSCPTNsGEDKQxNXta0U/8eJj/yZcig9wbmudYkl+MkdEoNTgsF24o
z+MOQld6XdLPythV4oX4FsRRkNl3Q4UVa7nWW1eu4I9fv+8uyw3usoD81kagzOmW
o0X6CgHbEsRORvzovDT3c8jxEafBH3+ou2mJ6Zv3gj8whbDx9+O8anHBmUs43Kwd
0e15IALgBo26K6xUnbQrL4vFHz+5G76SxYxpnhNgliGQUhG8ZRWedQ+MPrm6Ynja
CXG0LPb5ngWBn3/w3nqhHMl18DF74K5ldFUAL7r8hLvv0t2sqUa7AQrqDPHb/us3
4wJR3cOv4O25ryZdWU7vyDq9C9pnx2M1onQcY3W752g0Qu/D66v5H0CHuBMXyFu3
+mQ+K6taZYHEmZ5x7AOXcyC7Qx/qVhiPqNBCtEzbzmgtF7KqXyzbN+2cTDEInlIz
jLKMoZ1J8sNbhRmDqqqKhLq90NOQWz5wfDVHgD71SW2QRWbWZW+tMJqPwzp/b8kX
XxrUV/9J6MGlMhyl1dSOCn0bJ8zwyfiYeGLlUZ/pXv/vQaEqGDQqCmd0OJFzug+0
zh92RzCHGX/oE3tbeUoGQ/5S24jRMNS/oO8hBnx+vK1d2FPfj+w5N48ZsvrmEtpJ
dVlAE4KI8o7UIB1i4KaCHNb5Ae41VphhSy7k8icZELPRiuSfaGohRAVgAX7lB2iR
UXfCjwQFTFFGwmrokVLauWUEEDNzo6ZA7zHQJ79sL1GMaj9cQAZW0ktQ3t8agOq1
jhaKsHgVlvDtgsxkd8Zs1v78lRsCjjoXfqbeOgfFgh28Jd5nbeTgPusFbsk4iiAy
o5wAQgqqyg0NMRLNEnRa4l9QKQmD2fvtYU87OXSBJNmpv0vbCVNX8/6earR3JNvh
DAROLcpgCM6yCrV/lueZKQJ6EZd3acfqUKBgDC9vp9wBA25xBmOVd/M/MVOTa6Fn
5/44Xd2smABwZ5QduyihDKuyij9cch0bd7ThFbX5c7wWAAoGPIZ+yKcmDjG70cl9
HMV/5IF9qkcjoBkDAUw/e4NvG71OIk5Vl76Zh8dp0+An94H659VTq1d0gte9VgC2
kJz+fwHtpM0b7G1G5lCnV6sCJdlJgYZeZEk4sjTYegeEpuR7gCLmkBvXHcK76pvp
DQ7h2Wf6XvOzWQ7f80oNeOsj6y1boYM2m98JCZSb5zgyLVJ6xz5XvEJlTxHkBAbm
cohQ/NLDcXk3WY+BaD0j3HtECQWr8Pi/Y6fgv2mU5EH0kKk2i4XJzR1CBmVZKEjM
lBHAGD4QrTPYXEOmqWYYs5eCXAfeZNcBTF7d8lFGSsJwV0REwebjJHfe3E5DZock
vBuPjnY9gtA9Q6+JGluOocYL65NwUyRCwIKGrkL17/cc04K9otZXuD5noBRsXrq1
L8sfJ7kth1GMmNBwFR/Q4nPPALehjqp+6lOcHuM//Xn+Ll3WleSoD2JNi5BiaCTg
llUDYsgQUDKOdGOhBZd3c8z1mX451ceWAO5+7NZZttMras9is37vgLu2OHDlFWYm
g0xRzCv9UPqb0iKbbFonrlBCbiURRKiSgCSQ9spg03jewIqSqoxuJlJV1npzm64i
d6g7qN+xbB3+mRFT/zInj7X5maO0hN23Gakqdsb+AHFWwJJdv0Oi4E2R7zOTUP51
2JzKCyKolHi9fbx/wgarZWJojhdlVetHqC4sMKJWN8a3z3sS90MUWs5u+4i61cZK
hbbSN343gsHrldD9cP29Z9nzP8PWCLAWzT2DnDWH9vQQDJFqAyWTHCXLKpyIyUIx
1RbcOQ2nZup2P2SCoKzjlW3bGfQy+M9FlPDNx1u77jdWnr71W1NUuQwoq2Z9/C0Z
mLtAkUGm7/y4qeChifwDBuAQHmNVaWeFsac5DLlyCf/lTIkJiaEvQUMNPowXoh6f
ibBDxE214sRpNlXvh7R63SdvtOcQ0KgyKkcq1cdhcYaP0mKsGFgJ49bXKLA9yvJ+
bU4KSN2LugejpmOAwoxmHM+byLvMiBdeiMG1buhAcWyGXhyteGpbC3AB1GNUQVIu
0cb5G3RKdsjeOAn0twyksYNg0Yt9RvRDprG9TDNnqFSZk+w/xbEUjznPzXi7uOQ7
H/JDGLprJVSfoRXIPpT7Y2bGWkT4cFwIkBMsIU8nMr3ifd762KpKiPhgxiFcIw/t
6V11a5n3SE5TSMMpMIYmEaNtOIVFvB6Dr8gJNu4vPlcYHKOB5Kl+WB+CpBPAVIJA
/hml/qdnRKBtbkcvMCfiSdsH6QeZXn/zNGWA8uSXrVHFsBAGaByK2WDuOT36dtN2
t+t7+grmWe50O25c1H/RoT5y7KpfiogVZNZbTrXYDi8x4BNa5AkikApYCjhD820H
AKRM8qk1uCe89DyEVkkAEU8gkD3/y0MIjXnu+VyMfGsstIppRdcQsK+/rjKqHG3V
IpcdqpKxxfWkCMBsHhI/dSEAZY7Zvl4qJpfbC/u4J7BZGOR/GUzi5XqVAYd/LCJJ
2qMfFNpqV3SGC7A2cRZXjz/2QidqPuxpRlgZauSKYoniBl/DEp7hXCS2721X8xFp
5QVzjxgp4wU+j5bUnewgFY9ZJASpUD3e6n12+HhETYH8Xm7iVv+/5zasGsX1Yfal
HmaepoxPvN0OTkBxpz7pDLh7anUTUiq5y4E5pPbiH27mvFY+pV1afnH2F4bj4+lC
cNxHJ/ZBp/LJw9GphvMcUWZWKUUe/min8W8ZoLorRWJetIRnlT1qldD4TDrFH3B+
ckAb7Jxpaq0dKrIrcMWdbNbwfrl078BJBszU4zSJh1+D3uZDMJd/JLmmxECe04ll
cmCcgymo6JAwvqk3pF23+EnOmNofraEf6jgVRRoV0cPA9mgXXuLVFvUqKqBrFdY8
jLS8QghzxH72XC2pcSKFTS0FhmUmAy0kLsfoJ0aXvt9cdLqIJf90II3a39Kw0J1+
VRUASaFXr6Sd+mVGrMgYKJiXeVJMLaZcrvXOtt3VKeugosZ3l5MiWUQCVm3AnBhT
mt/PmqUbpEtUkmviCaMFmpCTms+uGQCIUvTmnRoZkfZ1Hdv8p45PYzRQ9Pdrb9Ox
zlGjndeeL8ufbJj/WrfZaOKNK27WK8o3xLJE4GvWXRaQdkHAUOw/lBU924ejhR7D
el7T/Y6BeskEFfa4u3VMF9yUsYYIlp4db9q9sQcjK+j3jrpGAZGlL6QS8mzQW8ji
9aHIQXKrrV4XnQlG0RaQfqKc8gcxQCDb4LhZ468PXjJQUY8lKPNv9aNkkOqw5pBK
cGB69ncyKIenTscJw7QFxo2Kw5Ayt/Y+y4JhGOZPGRPPmdc7Y+ghPqDgDDfIDysR
jy1n+JEVyF0ar8A1Dc3rRJfmEj4BeX9prORZXjd7rTqDZRwSB27c9dpMJE/Lklzn
SrUqt2q/MvcyWUbFBKklonFa+KA0xBILt/Fo1e1ad4KGjViwWE2yY9UqJsBofOOJ
UrT2Dyj8eMTJj8/1rd/tXFj/i4JV+NoNGd5pAfG45SbPMqaYJ+Kh/d+mYWWjCvaT
TmfZyXjmyzVW6pxGNUMaLZlTOO1IAiQCwLPD2eEVF1unTA2zcVjXpdkCoPbCgO7p
F9uiM3T4gbVBKy13egfApbiA/v7CH7BdAJS0rk+0nT212rQr2jEGYj0Tbm1bm0uf
cK2MsFrFoVy+BiPHOgsl7Dyb0mbFrK/fLEQ7TD7yd4Qq4UeMa8E0lz06RH0aQVXc
caToGmFgysFe0BS0Ck/64uLnllSuPPEoxba7tHyThIoDPcWOyOBRhADuuOAf7gNX
+L1lP0FCUucpd6Kyjrr1plmyCpiDYuMu7JOdALD0r5WOEeMQFwNiB9IEo63d8bax
I2K6FyD5OEdQEpwkWwc5KcFKtSVr1D3D8MDttFE7mnVnuh7JaI58cgkgRYIXX3pc
5/oTuu1VpEbxMtAHa2NPyGx/G5eoRsO/Lfohm0k9+DufBST0ZphIVKDATEATdy7y
F7NVoOCqKd3bsuui0NqIbfMtnhYInDDSwwwNJoPra5MrIZgxR3qu1bwToUrBBrlj
LDoEmgsbxM3cJaPm9++ZKPsIxifOlBxol/S63JjHYyl0kYjVihtGOPCG0hnGNz12
zZQXHB7a8TJojRGupoKmHXWI7gATEKygqOFrOFsu09l7M1yGLH7Ljo5FED8CE+mx
3Xex8aYhmR6zt+V0YtcNRzTWtMXPxMQ3yv6drDEm9ahWfmOLBvMXEiUedi8Q+L/e
kt4+2D0ARJylAO7nOWDX1lWYZS0s1NnfzQ+UE7GBswsKqJe2MzbazAYzr43yflsK
goPC2XDXJ1IkIX/enxRKFe7pTFhmCGroZExyH3f17PVjo0HWVvrJE1mATQPQvUaB
PluR4ZhWQfrXUoFvpB7/F0LF3CcAtmkpc4d5kiwee+KNZ0L/lo6VviEut5O4NyGB
2b9NYCznePtlKIVwbro1PR3eKKMWC2NUdDfqtZZRx5gKVwe/Z5obY4VT48qHlgUg
NHcerb9JlbdxWoaw6IafyjadHskosL8F1i1KgyeJ/Ci6SPiJdS9kYbcHaX7lDSN8
46QYAoRPmAdoUyTZbG6nxRtnqgWr41NrlyU0lWBRtaFyd3oXTWoSgIAf50o/6650
+OPah5+4Kq5isqLF/VdGQGD9aRjjSI1X4AW6k9/J0gdJHrZnwvMcdgVu91WVl5iE
+kcLKAeziFHWUBxsfdkjOV4J6Dm+PU1e8men3yjSVuS+BlQmKrBwAYzYejbvzTj7
IQAhOH4tqYn248kVDU/ANU5PtlAwBu/zwCeJmkU6zZLqgsmitJ4WopG+wx8SkrPq
V8zfzClyxVDlMBjYlIa8w4fz1GOOwTffgoFIBpdROLt4iB2iPJI/k+CXYYVmq+Q1
s2yw/sX6rRU78jLZpjLL+6O8yGR+SvBPDvpbQRomVB0mhC2BexcG8VLmlbbeCgLF
nyRYhbjezYmFUyrHUnbBZ/mh4/4A0b3rLcXgSwTZpNVWSk6ASneowEI4TgmdrCke
DKGr1R34duGbaEVFq+W5SfnegkH2KULsSloG8iHPsNmmfWrbXQabTbehW1RjSRHm
OFc/YnHa6f8ICpnS0QHEzaHf2q2osLPylNjviIdonWrzMzsObRSWLyb4xVb0LhEE
OlbADWE+lIgNLSymgQJGtCY5FnYYV8pZy4AgbTALf74myaLr7Lmuucw0A6GrWdgz
x8Uqc+ZwHYCj4K/uh7aSMspm+6lkyVvvMBFj6knk6TBXvoqWywE/m5w/iYp5LeZb
MD8jZMOHkCXfzwLDvXTpqEJJrLZiqgDU4pcJT+c/yH+9Dbp1g6FAkpLCzQPxaix5
KIVm4gzhnJspE3xUp/W7c+QEbKHbb4MavdHqrgHxdaMt2+38CTUvxXhKC20RXm/h
3hZui24Z8Ar8a55fdUX2VejbBrMi40afJBsg44fAEPcpsyaUjMq2eOmMn0cyj7Hf
UmUjCftwdpqga9WKqC7NSQp3/lspQ8X6+R2xjQjWGJg5g2LOpAz/eGF26LV67R4w
Wh033cks9zI+oXL3CJhCZwT3RwqJ8Dy+GbfteMadkRarHP1NvARgZmzJ1rYs8Hv8
k2fyb/UgwzAoBrOc50LUstpbo6vTTIWRrxYakCw2y5x5Kg1XiBGk6i3gwuEuhwB/
MNTa16CVIc4Jd6x0KbMoQVxdvlTF38kAq2572UO5rw7VpO02Yg1hnZewLdEHObbB
xtCLtrzWwdsrov7U8xskQDxgeS/gzc/trKAd90Na7BoctxLytiCJ9jq4EnwRgDIB
bzYG3GyS47CRtq5Fb/+MQDZW44W/wkWoqoKPYnpe9lI413KLa59srlPHFejJxZVE
JYRKJoKuCcSEV50MdKyIDqkMQAoFi2aurN8WlutCdZc6JEyadM/80dyDUaGGaUZB
Hob19YjuAW8kqFl+gAhxg9pI9xG3k3npOOqC6FD5pf0S4OhaW/aCa8tJX8R9+eZH
FcqLkNWIcxBKdpIlW24qgdoYIhxbr2TpOHr1Weswzt4nApGOgSJ85AdFGUObRth5
YXbq0KrqFruYMD+hbj3s1EHYXGQx/2k3mDw/YVgsOhFuaDFYfBbpnFgW1Hmg07jg
uvzyVFWJgJpSDPypFcHjqIuL5yaVvChaCspEl4C6WMD4nF7tiJMz6tytt8D8h6QO
iIAjGPPFEkMjJfeTNnLQAc3x9A/THE9tx2e4+o96LK4iel4JtLqJFG3uv5pjt7WW
JoYxd2dfPtVf2ZcQ639QqTSSycIimP1HZs/I5a8YnkDjK7WBpzcpLK2SDzevNjjt
ZBq4mHkqUK5jR9JYquEtoKdknOZy/TKgywFflJwqupWjLcVsNmDOsj2IeJDISSXv
cSkgIGJnoybXpo69SFEp4v8vIJyTMyHGzNIF4Wq/v99YHnWNkQPe7+7c222Mp8KV
YLROm38C0ZtdM/9+15gasOQYbTLlIPUR49+E0wss6IqUX2RPdl49UnD+4/kqCvRj
j/L36bO4mIu88LoGnE6bG0lhD4gDJbKRl1BuEdCocymOTcmEVEMn9g+6MgNWJpuV
hAVvnxIAyJkBaAyrg3GhfCpi1EpxowgXtyVp37JGNLlznUrgqBtZAEXNrBou06o5
+tqI0sXVm67xTSayNF0hb8npE4Rte3r8uu0OG/AyTbDiPPR0PZXm5xjlSUEYzcqK
lqYCbXSK4K7AA2Yn4LwjNba9Y4/aup5EPyx8/xaBNIz0vQ+TKQHyFI/gw52cvZ+c
h2ONQuHNGISuoVczAiwrHApzEv0972DW1w0x4KAu1SGj8mNMEP4b/TuKeIM4PMJW
/XmrjcszJt66TBG2dClBO/zIgVylLbJIIIcM1fxl1DtxBuwLDY9QdfuLRdqs4LI5
vtGRU1r+zD9qyMUOa5w4JvxfwKe1uKuYGE64gQtHiuaObjMV8qwLazC4Cbb01JwT
bn08ONN9amsAz1JzabiXCn+1p2KEe7Q8eCHvjkYmrMKuG5D6Wyy+yjCTndA2rxZB
iqFbmFDlKeIrJh1xMQ/xn0hksG1MoApJM+l+JAMH+/dIc1+vjvjluvjPpBPz21gA
u9YihTe4WFqHE9VZoDmHHS/u9zItG31o19hDnGJcH9XU9x0B1kfKYcdUwchYDWyP
qpFzSJrEEMlUZ6gtyLF9KZSi4QTukPqwSlqlfj+6K8lY1oOZ1+fVC32/unRWuH6O
Ud+HzirJ98sFiaykY27vMqEBB2lFEbY6TA6jd/96j8oVJi45zE266Iiwe7VjVszD
1XXjYakzxVNYWZDFUEs6BRKD6MU89IxNtjZOK7boWoHb14P9Azse1CufX1MDZhK2
2hxSkbudnIdlj8nUv5yQyCL0uX1ujZjvKywkdmFpTIQtZNY4itVHK4q9/tvzufBG
fPyF9Fe2cA5OqLOhopx0VIRghd+ddlb6/xKBS/52snJv+h0HcT1HVJ7OyZeaL3us
1xfxKu8leu8dX5Fyyg3W963ZluKCPhbhf2cie3j0xPzE2Fc2Nq+aX2AONzM6MwzP
WPc0NtZk1RE90UqSqyZ9ZwPQg9k738aL6WBDXj/v3YtbCkKNdxUSOtim2qyRuUiX
//pragma protect end_data_block
//pragma protect digest_block
hj8PnBEKKogeOKVu0W8h1SB9q8w=
//pragma protect end_digest_block
//pragma protect end_protected
